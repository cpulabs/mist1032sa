/*****************************************************************************************************
Files that are included in this project is deliverable by all Open Design Computer Project.
http://open-arch.org

All files included in this project have been allocated in the BSD licence.	
Open Design Computer Project @Takahiro Ito
	
Make	:	2012/08/04
*****************************************************************************************************/

`default_nettype none


`define		LOAD_WORD			32'd10000//32'd1024
`define		WAIT_CYCLE			32'd1200//32'h2028



module debug_rom(
				//System
				input				iCLOCK,
				input				inRESET,
				//Debugg
				output				oDEBUG_VALID,
				output				oDEBUG_MEMIF_REQ_VALID,
				output				oDEBUG_MEMIF_REQ_DQM0,
				output				oDEBUG_MEMIF_REQ_DQM1,
				output				oDEBUG_MEMIF_REQ_DQM2,
				output				oDEBUG_MEMIF_REQ_DQM3,
				output				oDEBUG_MEMIF_REQ_RW,
				output	[24:0]		oDEBUG_MEMIF_REQ_ADDR,
				output	[31:0]		oDEBUG_MEMIF_REQ_DATA,
				input				iDEBUG_MEMIF_REQ_LOCK
	);
		
	//END Controll
	reg					b_write_end;
	reg					b_wait_end;
	reg		[31:0]		b_write_counter;
	reg		[31:0]		b_wait_counter;
	always@(posedge iCLOCK or negedge inRESET)begin
		if(!inRESET)begin
			b_write_end			<=		1'b0;
			b_wait_end			<=		1'b0;
			b_write_counter		<=		32'h0;
			b_wait_counter		<=		32'h0;
		end
		else begin
			if(!b_write_end)begin
				if(!iDEBUG_MEMIF_REQ_LOCK)begin
					b_write_counter		<=		b_write_counter + 32'h1;
				end
				if(b_write_counter == `LOAD_WORD)begin
					b_write_end			<=		1'b1;
				end
			end
			else begin
				b_write_end			<=		1'b1;
				if(!b_wait_end)begin
					b_wait_counter		<=		b_wait_counter + 32'h1;
					if(b_wait_counter == `WAIT_CYCLE)begin
						b_wait_end			<=		1'b1;
					end
				end
			end
		end
	end
	
	
	

	
	function [31:0] func_rom_io_display_test;
		input	[31:0]		func_addr;
		begin
			case(func_addr)	
				//Dhrystone
				0		:	func_rom_io_display_test	=	32'h0ee08000;		//[0]lih      r0,0x400
				1		:	func_rom_io_display_test	=	32'h1c000000;		//[4]srspw    r0
				2		:	func_rom_io_display_test	=	32'h110003e0;		//[8]push     rret
				3		:	func_rom_io_display_test	=	32'h207003e2;		//[C]movepc   rret,8
				4		:	func_rom_io_display_test	=	32'h143000f4;		//[10]br       3e0 <start>,#al
				5		:	func_rom_io_display_test	=	32'h14300000;		//[14]br       14 <_start+0x14>,#al
				8		:	func_rom_io_display_test	=	32'h110003c0;		//[20]push     rbase
				9		:	func_rom_io_display_test	=	32'h180003c0;		//[24]srspr    rbase
				10		:	func_rom_io_display_test	=	32'h0ee00040;		//[28]lih      r2,0x0
				11		:	func_rom_io_display_test	=	32'h0d498450;		//[2C]wl16     r2,0x4c30
				12		:	func_rom_io_display_test	=	32'h10400002;		//[30]ld32     r0,r2
				13		:	func_rom_io_display_test	=	32'h00200001;		//[34]sub      r0,r1
				14		:	func_rom_io_display_test	=	32'h0edffc3c;		//[38]lil      r1,-4
				15		:	func_rom_io_display_test	=	32'h0c000001;		//[3C]and      r0,r1
				16		:	func_rom_io_display_test	=	32'h10a00002;		//[40]st32     r0,r2
				17		:	func_rom_io_display_test	=	32'h120003c0;		//[44]pop      rbase
				18		:	func_rom_io_display_test	=	32'h144003e0;		//[48]b        rret,#al
				19		:	func_rom_io_display_test	=	32'h00000000;		//[4C]add      r0,r0
				20		:	func_rom_io_display_test	=	32'h110003c0;		//[50]push     rbase
				21		:	func_rom_io_display_test	=	32'h180003c0;		//[54]srspr    rbase
				22		:	func_rom_io_display_test	=	32'h10400061;		//[58]ld32     r3,r1
				23		:	func_rom_io_display_test	=	32'h0ee00000;		//[5C]lih      r0,0x0
				24		:	func_rom_io_display_test	=	32'h0d4e6c0c;		//[60]wl16     r0,0x736c
				25		:	func_rom_io_display_test	=	32'h10000000;		//[64]ld8      r0,r0
				26		:	func_rom_io_display_test	=	32'h03800040;		//[68]sext8    r2,r0
				27		:	func_rom_io_display_test	=	32'h00d00841;		//[6C]cmp      r2,65
				28		:	func_rom_io_display_test	=	32'h14320008;		//[70]br       90 <Proc_2+0x40>,#neq
				29		:	func_rom_io_display_test	=	32'h20400003;		//[74]move     r0,r3
				30		:	func_rom_io_display_test	=	32'h00100009;		//[78]add      r0,9
				31		:	func_rom_io_display_test	=	32'h0ee00040;		//[7C]lih      r2,0x0
				32		:	func_rom_io_display_test	=	32'h0d4e6c48;		//[80]wl16     r2,0x7368
				33		:	func_rom_io_display_test	=	32'h10400042;		//[84]ld32     r2,r2
				34		:	func_rom_io_display_test	=	32'h00200002;		//[88]sub      r0,r2
				35		:	func_rom_io_display_test	=	32'h10a00001;		//[8C]st32     r0,r1
				36		:	func_rom_io_display_test	=	32'h120003c0;		//[90]pop      rbase
				37		:	func_rom_io_display_test	=	32'h144003e0;		//[94]b        rret,#al
				40		:	func_rom_io_display_test	=	32'h110003c0;		//[A0]push     rbase
				41		:	func_rom_io_display_test	=	32'h110003e0;		//[A4]push     rret
				42		:	func_rom_io_display_test	=	32'h180003c0;		//[A8]srspr    rbase
				43		:	func_rom_io_display_test	=	32'h0ee00060;		//[AC]lih      r3,0x0
				44		:	func_rom_io_display_test	=	32'h0d4e6c70;		//[B0]wl16     r3,0x7370
				45		:	func_rom_io_display_test	=	32'h10400003;		//[B4]ld32     r0,r3
				46		:	func_rom_io_display_test	=	32'h00d00000;		//[B8]cmp      r0,0
				47		:	func_rom_io_display_test	=	32'h14310010;		//[BC]br       fc <Proc_3+0x5c>,#eq
				48		:	func_rom_io_display_test	=	32'h10400000;		//[C0]ld32     r0,r0
				49		:	func_rom_io_display_test	=	32'h10a00001;		//[C4]st32     r0,r1
				50		:	func_rom_io_display_test	=	32'h10400063;		//[C8]ld32     r3,r3
				51		:	func_rom_io_display_test	=	32'h0ee00040;		//[CC]lih      r2,0x0
				52		:	func_rom_io_display_test	=	32'h0d4e6c48;		//[D0]wl16     r2,0x7368
				53		:	func_rom_io_display_test	=	32'h0ec0002a;		//[D4]lil      r1,10
				54		:	func_rom_io_display_test	=	32'h10400042;		//[D8]ld32     r2,r2
				55		:	func_rom_io_display_test	=	32'h0010006c;		//[DC]add      r3,12
				56		:	func_rom_io_display_test	=	32'h0ee003a0;		//[E0]lih      rtmp,0x0
				57		:	func_rom_io_display_test	=	32'h0d411fb0;		//[E4]wl16     rtmp,0x8f0
				58		:	func_rom_io_display_test	=	32'h207003e2;		//[E8]movepc   rret,8
				59		:	func_rom_io_display_test	=	32'h144003a0;		//[EC]b        rtmp,#al
				60		:	func_rom_io_display_test	=	32'h120003e0;		//[F0]pop      rret
				61		:	func_rom_io_display_test	=	32'h120003c0;		//[F4]pop      rbase
				62		:	func_rom_io_display_test	=	32'h144003e0;		//[F8]b        rret,#al
				63		:	func_rom_io_display_test	=	32'h20400060;		//[FC]move     r3,r0
				64		:	func_rom_io_display_test	=	32'h1430fff3;		//[100]br       cc <Proc_3+0x2c>,#al
				68		:	func_rom_io_display_test	=	32'h110003c0;		//[110]push     rbase
				69		:	func_rom_io_display_test	=	32'h11000200;		//[114]push     r16
				70		:	func_rom_io_display_test	=	32'h11000220;		//[118]push     r17
				71		:	func_rom_io_display_test	=	32'h11000240;		//[11C]push     r18
				72		:	func_rom_io_display_test	=	32'h11000260;		//[120]push     r19
				73		:	func_rom_io_display_test	=	32'h11000280;		//[124]push     r20
				74		:	func_rom_io_display_test	=	32'h110002a0;		//[128]push     r21
				75		:	func_rom_io_display_test	=	32'h110002c0;		//[12C]push     r22
				76		:	func_rom_io_display_test	=	32'h110003e0;		//[130]push     rret
				77		:	func_rom_io_display_test	=	32'h180003c0;		//[134]srspr    rbase
				78		:	func_rom_io_display_test	=	32'h20400221;		//[138]move     r17,r1
				79		:	func_rom_io_display_test	=	32'h10400201;		//[13C]ld32     r16,r1
				80		:	func_rom_io_display_test	=	32'h0ee00240;		//[140]lih      r18,0x0
				81		:	func_rom_io_display_test	=	32'h0d4e6e50;		//[144]wl16     r18,0x7370
				82		:	func_rom_io_display_test	=	32'h10400012;		//[148]ld32     r0,r18
				83		:	func_rom_io_display_test	=	32'h10400020;		//[14C]ld32     r1,r0
				84		:	func_rom_io_display_test	=	32'h10a00030;		//[150]st32     r1,r16
				85		:	func_rom_io_display_test	=	32'h20400290;		//[154]move     r20,r16
				86		:	func_rom_io_display_test	=	32'h00100284;		//[158]add      r20,4
				87		:	func_rom_io_display_test	=	32'h20400020;		//[15C]move     r1,r0
				88		:	func_rom_io_display_test	=	32'h00100024;		//[160]add      r1,4
				89		:	func_rom_io_display_test	=	32'h10400021;		//[164]ld32     r1,r1
				90		:	func_rom_io_display_test	=	32'h10a00034;		//[168]st32     r1,r20
				91		:	func_rom_io_display_test	=	32'h204002d0;		//[16C]move     r22,r16
				92		:	func_rom_io_display_test	=	32'h001002c8;		//[170]add      r22,8
				93		:	func_rom_io_display_test	=	32'h20400020;		//[174]move     r1,r0
				94		:	func_rom_io_display_test	=	32'h00100028;		//[178]add      r1,8
				95		:	func_rom_io_display_test	=	32'h10400021;		//[17C]ld32     r1,r1
				96		:	func_rom_io_display_test	=	32'h10a00036;		//[180]st32     r1,r22
				97		:	func_rom_io_display_test	=	32'h20400270;		//[184]move     r19,r16
				98		:	func_rom_io_display_test	=	32'h0010026c;		//[188]add      r19,12
				99		:	func_rom_io_display_test	=	32'h20400020;		//[18C]move     r1,r0
				100		:	func_rom_io_display_test	=	32'h0010002c;		//[190]add      r1,12
				101		:	func_rom_io_display_test	=	32'h10400021;		//[194]ld32     r1,r1
				102		:	func_rom_io_display_test	=	32'h10a00033;		//[198]st32     r1,r19
				103		:	func_rom_io_display_test	=	32'h20400050;		//[19C]move     r2,r16
				104		:	func_rom_io_display_test	=	32'h00100050;		//[1A0]add      r2,16
				105		:	func_rom_io_display_test	=	32'h20400020;		//[1A4]move     r1,r0
				106		:	func_rom_io_display_test	=	32'h00100030;		//[1A8]add      r1,16
				107		:	func_rom_io_display_test	=	32'h10400021;		//[1AC]ld32     r1,r1
				108		:	func_rom_io_display_test	=	32'h10a00022;		//[1B0]st32     r1,r2
				109		:	func_rom_io_display_test	=	32'h00100044;		//[1B4]add      r2,4
				110		:	func_rom_io_display_test	=	32'h20400020;		//[1B8]move     r1,r0
				111		:	func_rom_io_display_test	=	32'h00100034;		//[1BC]add      r1,20
				112		:	func_rom_io_display_test	=	32'h10400021;		//[1C0]ld32     r1,r1
				113		:	func_rom_io_display_test	=	32'h10a00022;		//[1C4]st32     r1,r2
				114		:	func_rom_io_display_test	=	32'h00100044;		//[1C8]add      r2,4
				115		:	func_rom_io_display_test	=	32'h20400020;		//[1CC]move     r1,r0
				116		:	func_rom_io_display_test	=	32'h00100038;		//[1D0]add      r1,24
				117		:	func_rom_io_display_test	=	32'h10400021;		//[1D4]ld32     r1,r1
				118		:	func_rom_io_display_test	=	32'h10a00022;		//[1D8]st32     r1,r2
				119		:	func_rom_io_display_test	=	32'h00100044;		//[1DC]add      r2,4
				120		:	func_rom_io_display_test	=	32'h20400020;		//[1E0]move     r1,r0
				121		:	func_rom_io_display_test	=	32'h0010003c;		//[1E4]add      r1,28
				122		:	func_rom_io_display_test	=	32'h10400021;		//[1E8]ld32     r1,r1
				123		:	func_rom_io_display_test	=	32'h10a00022;		//[1EC]st32     r1,r2
				124		:	func_rom_io_display_test	=	32'h00100044;		//[1F0]add      r2,4
				125		:	func_rom_io_display_test	=	32'h20400020;		//[1F4]move     r1,r0
				126		:	func_rom_io_display_test	=	32'h00100420;		//[1F8]add      r1,32
				127		:	func_rom_io_display_test	=	32'h10400021;		//[1FC]ld32     r1,r1
				128		:	func_rom_io_display_test	=	32'h10a00022;		//[200]st32     r1,r2
				129		:	func_rom_io_display_test	=	32'h00100044;		//[204]add      r2,4
				130		:	func_rom_io_display_test	=	32'h20400020;		//[208]move     r1,r0
				131		:	func_rom_io_display_test	=	32'h00100424;		//[20C]add      r1,36
				132		:	func_rom_io_display_test	=	32'h10400021;		//[210]ld32     r1,r1
				133		:	func_rom_io_display_test	=	32'h10a00022;		//[214]st32     r1,r2
				134		:	func_rom_io_display_test	=	32'h00100044;		//[218]add      r2,4
				135		:	func_rom_io_display_test	=	32'h20400020;		//[21C]move     r1,r0
				136		:	func_rom_io_display_test	=	32'h00100428;		//[220]add      r1,40
				137		:	func_rom_io_display_test	=	32'h10400021;		//[224]ld32     r1,r1
				138		:	func_rom_io_display_test	=	32'h10a00022;		//[228]st32     r1,r2
				139		:	func_rom_io_display_test	=	32'h20400030;		//[22C]move     r1,r16
				140		:	func_rom_io_display_test	=	32'h0010042c;		//[230]add      r1,44
				141		:	func_rom_io_display_test	=	32'h0010040c;		//[234]add      r0,44
				142		:	func_rom_io_display_test	=	32'h10400000;		//[238]ld32     r0,r0
				143		:	func_rom_io_display_test	=	32'h10a00001;		//[23C]st32     r0,r1
				144		:	func_rom_io_display_test	=	32'h204002b1;		//[240]move     r21,r17
				145		:	func_rom_io_display_test	=	32'h001002ac;		//[244]add      r21,12
				146		:	func_rom_io_display_test	=	32'h0ec00005;		//[248]lil      r0,5
				147		:	func_rom_io_display_test	=	32'h10a00015;		//[24C]st32     r0,r21
				148		:	func_rom_io_display_test	=	32'h10a00013;		//[250]st32     r0,r19
				149		:	func_rom_io_display_test	=	32'h10400011;		//[254]ld32     r0,r17
				150		:	func_rom_io_display_test	=	32'h10a00010;		//[258]st32     r0,r16
				151		:	func_rom_io_display_test	=	32'h20400030;		//[25C]move     r1,r16
				152		:	func_rom_io_display_test	=	32'h0ee003a0;		//[260]lih      rtmp,0x0
				153		:	func_rom_io_display_test	=	32'h0d4017a0;		//[264]wl16     rtmp,0xa0
				154		:	func_rom_io_display_test	=	32'h207003e2;		//[268]movepc   rret,8
				155		:	func_rom_io_display_test	=	32'h144003a0;		//[26C]b        rtmp,#al
				156		:	func_rom_io_display_test	=	32'h10400294;		//[270]ld32     r20,r20
				157		:	func_rom_io_display_test	=	32'h00d00280;		//[274]cmp      r20,0
				158		:	func_rom_io_display_test	=	32'h14310044;		//[278]br       388 <Proc_1+0x278>,#eq
				159		:	func_rom_io_display_test	=	32'h10400011;		//[27C]ld32     r0,r17
				160		:	func_rom_io_display_test	=	32'h10400020;		//[280]ld32     r1,r0
				161		:	func_rom_io_display_test	=	32'h10a00031;		//[284]st32     r1,r17
				162		:	func_rom_io_display_test	=	32'h20400051;		//[288]move     r2,r17
				163		:	func_rom_io_display_test	=	32'h00100044;		//[28C]add      r2,4
				164		:	func_rom_io_display_test	=	32'h20400020;		//[290]move     r1,r0
				165		:	func_rom_io_display_test	=	32'h00100024;		//[294]add      r1,4
				166		:	func_rom_io_display_test	=	32'h10400021;		//[298]ld32     r1,r1
				167		:	func_rom_io_display_test	=	32'h10a00022;		//[29C]st32     r1,r2
				168		:	func_rom_io_display_test	=	32'h00100044;		//[2A0]add      r2,4
				169		:	func_rom_io_display_test	=	32'h20400020;		//[2A4]move     r1,r0
				170		:	func_rom_io_display_test	=	32'h00100028;		//[2A8]add      r1,8
				171		:	func_rom_io_display_test	=	32'h10400021;		//[2AC]ld32     r1,r1
				172		:	func_rom_io_display_test	=	32'h10a00022;		//[2B0]st32     r1,r2
				173		:	func_rom_io_display_test	=	32'h20400020;		//[2B4]move     r1,r0
				174		:	func_rom_io_display_test	=	32'h0010002c;		//[2B8]add      r1,12
				175		:	func_rom_io_display_test	=	32'h10400021;		//[2BC]ld32     r1,r1
				176		:	func_rom_io_display_test	=	32'h10a00035;		//[2C0]st32     r1,r21
				177		:	func_rom_io_display_test	=	32'h00100048;		//[2C4]add      r2,8
				178		:	func_rom_io_display_test	=	32'h20400020;		//[2C8]move     r1,r0
				179		:	func_rom_io_display_test	=	32'h00100030;		//[2CC]add      r1,16
				180		:	func_rom_io_display_test	=	32'h10400021;		//[2D0]ld32     r1,r1
				181		:	func_rom_io_display_test	=	32'h10a00022;		//[2D4]st32     r1,r2
				182		:	func_rom_io_display_test	=	32'h00100044;		//[2D8]add      r2,4
				183		:	func_rom_io_display_test	=	32'h20400020;		//[2DC]move     r1,r0
				184		:	func_rom_io_display_test	=	32'h00100034;		//[2E0]add      r1,20
				185		:	func_rom_io_display_test	=	32'h10400021;		//[2E4]ld32     r1,r1
				186		:	func_rom_io_display_test	=	32'h10a00022;		//[2E8]st32     r1,r2
				187		:	func_rom_io_display_test	=	32'h00100044;		//[2EC]add      r2,4
				188		:	func_rom_io_display_test	=	32'h20400020;		//[2F0]move     r1,r0
				189		:	func_rom_io_display_test	=	32'h00100038;		//[2F4]add      r1,24
				190		:	func_rom_io_display_test	=	32'h10400021;		//[2F8]ld32     r1,r1
				191		:	func_rom_io_display_test	=	32'h10a00022;		//[2FC]st32     r1,r2
				192		:	func_rom_io_display_test	=	32'h00100044;		//[300]add      r2,4
				193		:	func_rom_io_display_test	=	32'h20400020;		//[304]move     r1,r0
				194		:	func_rom_io_display_test	=	32'h0010003c;		//[308]add      r1,28
				195		:	func_rom_io_display_test	=	32'h10400021;		//[30C]ld32     r1,r1
				196		:	func_rom_io_display_test	=	32'h10a00022;		//[310]st32     r1,r2
				197		:	func_rom_io_display_test	=	32'h00100044;		//[314]add      r2,4
				198		:	func_rom_io_display_test	=	32'h20400020;		//[318]move     r1,r0
				199		:	func_rom_io_display_test	=	32'h00100420;		//[31C]add      r1,32
				200		:	func_rom_io_display_test	=	32'h10400021;		//[320]ld32     r1,r1
				201		:	func_rom_io_display_test	=	32'h10a00022;		//[324]st32     r1,r2
				202		:	func_rom_io_display_test	=	32'h00100044;		//[328]add      r2,4
				203		:	func_rom_io_display_test	=	32'h20400020;		//[32C]move     r1,r0
				204		:	func_rom_io_display_test	=	32'h00100424;		//[330]add      r1,36
				205		:	func_rom_io_display_test	=	32'h10400021;		//[334]ld32     r1,r1
				206		:	func_rom_io_display_test	=	32'h10a00022;		//[338]st32     r1,r2
				207		:	func_rom_io_display_test	=	32'h00100044;		//[33C]add      r2,4
				208		:	func_rom_io_display_test	=	32'h20400020;		//[340]move     r1,r0
				209		:	func_rom_io_display_test	=	32'h00100428;		//[344]add      r1,40
				210		:	func_rom_io_display_test	=	32'h10400021;		//[348]ld32     r1,r1
				211		:	func_rom_io_display_test	=	32'h10a00022;		//[34C]st32     r1,r2
				212		:	func_rom_io_display_test	=	32'h0010062c;		//[350]add      r17,44
				213		:	func_rom_io_display_test	=	32'h0010040c;		//[354]add      r0,44
				214		:	func_rom_io_display_test	=	32'h10400000;		//[358]ld32     r0,r0
				215		:	func_rom_io_display_test	=	32'h10a00011;		//[35C]st32     r0,r17
				216		:	func_rom_io_display_test	=	32'h120003e0;		//[360]pop      rret
				217		:	func_rom_io_display_test	=	32'h120002c0;		//[364]pop      r22
				218		:	func_rom_io_display_test	=	32'h120002a0;		//[368]pop      r21
				219		:	func_rom_io_display_test	=	32'h12000280;		//[36C]pop      r20
				220		:	func_rom_io_display_test	=	32'h12000260;		//[370]pop      r19
				221		:	func_rom_io_display_test	=	32'h12000240;		//[374]pop      r18
				222		:	func_rom_io_display_test	=	32'h12000220;		//[378]pop      r17
				223		:	func_rom_io_display_test	=	32'h12000200;		//[37C]pop      r16
				224		:	func_rom_io_display_test	=	32'h120003c0;		//[380]pop      rbase
				225		:	func_rom_io_display_test	=	32'h144003e0;		//[384]b        rret,#al
				226		:	func_rom_io_display_test	=	32'h0ec00006;		//[388]lil      r0,6
				227		:	func_rom_io_display_test	=	32'h10a00013;		//[38C]st32     r0,r19
				228		:	func_rom_io_display_test	=	32'h00100228;		//[390]add      r17,8
				229		:	func_rom_io_display_test	=	32'h10400031;		//[394]ld32     r1,r17
				230		:	func_rom_io_display_test	=	32'h20400056;		//[398]move     r2,r22
				231		:	func_rom_io_display_test	=	32'h0ee003a0;		//[39C]lih      rtmp,0x0
				232		:	func_rom_io_display_test	=	32'h0d410fa0;		//[3A0]wl16     rtmp,0x860
				233		:	func_rom_io_display_test	=	32'h207003e2;		//[3A4]movepc   rret,8
				234		:	func_rom_io_display_test	=	32'h144003a0;		//[3A8]b        rtmp,#al
				235		:	func_rom_io_display_test	=	32'h10400252;		//[3AC]ld32     r18,r18
				236		:	func_rom_io_display_test	=	32'h10400252;		//[3B0]ld32     r18,r18
				237		:	func_rom_io_display_test	=	32'h10a00250;		//[3B4]st32     r18,r16
				238		:	func_rom_io_display_test	=	32'h10400033;		//[3B8]ld32     r1,r19
				239		:	func_rom_io_display_test	=	32'h0ec0004a;		//[3BC]lil      r2,10
				240		:	func_rom_io_display_test	=	32'h20400073;		//[3C0]move     r3,r19
				241		:	func_rom_io_display_test	=	32'h0ee003a0;		//[3C4]lih      rtmp,0x0
				242		:	func_rom_io_display_test	=	32'h0d411fb0;		//[3C8]wl16     rtmp,0x8f0
				243		:	func_rom_io_display_test	=	32'h207003e2;		//[3CC]movepc   rret,8
				244		:	func_rom_io_display_test	=	32'h144003a0;		//[3D0]b        rtmp,#al
				245		:	func_rom_io_display_test	=	32'h1430ffe3;		//[3D4]br       360 <Proc_1+0x250>,#al
				248		:	func_rom_io_display_test	=	32'h110003c0;		//[3E0]push     rbase
				249		:	func_rom_io_display_test	=	32'h11000200;		//[3E4]push     r16
				250		:	func_rom_io_display_test	=	32'h11000220;		//[3E8]push     r17
				251		:	func_rom_io_display_test	=	32'h11000240;		//[3EC]push     r18
				252		:	func_rom_io_display_test	=	32'h11000260;		//[3F0]push     r19
				253		:	func_rom_io_display_test	=	32'h11000280;		//[3F4]push     r20
				254		:	func_rom_io_display_test	=	32'h110002a0;		//[3F8]push     r21
				255		:	func_rom_io_display_test	=	32'h110002c0;		//[3FC]push     r22
				256		:	func_rom_io_display_test	=	32'h110002e0;		//[400]push     r23
				257		:	func_rom_io_display_test	=	32'h11000300;		//[404]push     r24
				258		:	func_rom_io_display_test	=	32'h11000320;		//[408]push     r25
				259		:	func_rom_io_display_test	=	32'h11000340;		//[40C]push     r26
				260		:	func_rom_io_display_test	=	32'h11000360;		//[410]push     r27
				261		:	func_rom_io_display_test	=	32'h110003e0;		//[414]push     rret
				262		:	func_rom_io_display_test	=	32'h180003a0;		//[418]srspr    rtmp
				263		:	func_rom_io_display_test	=	32'h0010f7b4;		//[41C]add      rtmp,-76
				264		:	func_rom_io_display_test	=	32'h1c0003a0;		//[420]srspw    rtmp
				265		:	func_rom_io_display_test	=	32'h180003c0;		//[424]srspr    rbase
				266		:	func_rom_io_display_test	=	32'h0ee00040;		//[428]lih      r2,0x0
				267		:	func_rom_io_display_test	=	32'h0d498450;		//[42C]wl16     r2,0x4c30
				268		:	func_rom_io_display_test	=	32'h10400002;		//[430]ld32     r0,r2
				269		:	func_rom_io_display_test	=	32'h0ed80020;		//[434]lil      r1,-16384
				270		:	func_rom_io_display_test	=	32'h00000001;		//[438]add      r0,r1
				271		:	func_rom_io_display_test	=	32'h0edffc3c;		//[43C]lil      r1,-4
				272		:	func_rom_io_display_test	=	32'h0c000001;		//[440]and      r0,r1
				273		:	func_rom_io_display_test	=	32'h0010f810;		//[444]add      r0,-48
				274		:	func_rom_io_display_test	=	32'h0ee00020;		//[448]lih      r1,0x0
				275		:	func_rom_io_display_test	=	32'h0d4e6c24;		//[44C]wl16     r1,0x7364
				276		:	func_rom_io_display_test	=	32'h10a00001;		//[450]st32     r0,r1
				277		:	func_rom_io_display_test	=	32'h20400020;		//[454]move     r1,r0
				278		:	func_rom_io_display_test	=	32'h0010f830;		//[458]add      r1,-48
				279		:	func_rom_io_display_test	=	32'h10a00022;		//[45C]st32     r1,r2
				280		:	func_rom_io_display_test	=	32'h0ee00300;		//[460]lih      r24,0x0
				281		:	func_rom_io_display_test	=	32'h0d4e6f10;		//[464]wl16     r24,0x7370
				282		:	func_rom_io_display_test	=	32'h10a00038;		//[468]st32     r1,r24
				283		:	func_rom_io_display_test	=	32'h10a00001;		//[46C]st32     r0,r1
				284		:	func_rom_io_display_test	=	32'h0010f814;		//[470]add      r0,-44
				285		:	func_rom_io_display_test	=	32'h0ec00040;		//[474]lil      r2,0
				286		:	func_rom_io_display_test	=	32'h10a00040;		//[478]st32     r2,r0
				287		:	func_rom_io_display_test	=	32'h00100004;		//[47C]add      r0,4
				288		:	func_rom_io_display_test	=	32'h0ec00042;		//[480]lil      r2,2
				289		:	func_rom_io_display_test	=	32'h10a00040;		//[484]st32     r2,r0
				290		:	func_rom_io_display_test	=	32'h00100004;		//[488]add      r0,4
				291		:	func_rom_io_display_test	=	32'h0ec00448;		//[48C]lil      r2,40
				292		:	func_rom_io_display_test	=	32'h10a00040;		//[490]st32     r2,r0
				293		:	func_rom_io_display_test	=	32'h00100030;		//[494]add      r1,16
				294		:	func_rom_io_display_test	=	32'h0ee00040;		//[498]lih      r2,0x0
				295		:	func_rom_io_display_test	=	32'h0d417050;		//[49C]wl16     r2,0xb90
				296		:	func_rom_io_display_test	=	32'h0ee003a0;		//[4A0]lih      rtmp,0x0
				297		:	func_rom_io_display_test	=	32'h0d416bb0;		//[4A4]wl16     rtmp,0xb50
				298		:	func_rom_io_display_test	=	32'h207003e2;		//[4A8]movepc   rret,8
				299		:	func_rom_io_display_test	=	32'h144003a0;		//[4AC]b        rtmp,#al
				300		:	func_rom_io_display_test	=	32'h2040003e;		//[4B0]move     r1,rbase
				301		:	func_rom_io_display_test	=	32'h00100428;		//[4B4]add      r1,40
				302		:	func_rom_io_display_test	=	32'h0ee00040;		//[4B8]lih      r2,0x0
				303		:	func_rom_io_display_test	=	32'h0d417450;		//[4BC]wl16     r2,0xbb0
				304		:	func_rom_io_display_test	=	32'h0ee003a0;		//[4C0]lih      rtmp,0x0
				305		:	func_rom_io_display_test	=	32'h0d416bb0;		//[4C4]wl16     rtmp,0xb50
				306		:	func_rom_io_display_test	=	32'h207003e2;		//[4C8]movepc   rret,8
				307		:	func_rom_io_display_test	=	32'h144003a0;		//[4CC]b        rtmp,#al
				308		:	func_rom_io_display_test	=	32'h0ee00000;		//[4D0]lih      r0,0x0
				309		:	func_rom_io_display_test	=	32'h0d498810;		//[4D4]wl16     r0,0x4c50
				310		:	func_rom_io_display_test	=	32'h0ec0c85c;		//[4D8]lil      r2,1628
				311		:	func_rom_io_display_test	=	32'h00000002;		//[4DC]add      r0,r2
				312		:	func_rom_io_display_test	=	32'h0ec0002a;		//[4E0]lil      r1,10
				313		:	func_rom_io_display_test	=	32'h10a00020;		//[4E4]st32     r1,r0
				314		:	func_rom_io_display_test	=	32'h0ee003a0;		//[4E8]lih      rtmp,0x0
				315		:	func_rom_io_display_test	=	32'h0d415bb0;		//[4EC]wl16     rtmp,0xad0
				316		:	func_rom_io_display_test	=	32'h207003e2;		//[4F0]movepc   rret,8
				317		:	func_rom_io_display_test	=	32'h144003a0;		//[4F4]b        rtmp,#al
				318		:	func_rom_io_display_test	=	32'h0ee00040;		//[4F8]lih      r2,0x0
				319		:	func_rom_io_display_test	=	32'h0ec00828;		//[4FC]lil      r1,72
				320		:	func_rom_io_display_test	=	32'h0000003e;		//[500]add      r1,rbase
				321		:	func_rom_io_display_test	=	32'h0d498844;		//[504]wl16     r2,0x4c44
				322		:	func_rom_io_display_test	=	32'h10a00041;		//[508]st32     r2,r1
				323		:	func_rom_io_display_test	=	32'h10a00002;		//[50C]st32     r0,r2
				324		:	func_rom_io_display_test	=	32'h0ec00281;		//[510]lil      r20,1
				325		:	func_rom_io_display_test	=	32'h0ee00320;		//[514]lih      r25,0x0
				326		:	func_rom_io_display_test	=	32'h0d4e6f2c;		//[518]wl16     r25,0x736c
				327		:	func_rom_io_display_test	=	32'h0ee00260;		//[51C]lih      r19,0x0
				328		:	func_rom_io_display_test	=	32'h0d4e8a68;		//[520]wl16     r19,0x7448
				329		:	func_rom_io_display_test	=	32'h0ee00240;		//[524]lih      r18,0x0
				330		:	func_rom_io_display_test	=	32'h0d4e6e4d;		//[528]wl16     r18,0x736d
				331		:	func_rom_io_display_test	=	32'h204002de;		//[52C]move     r22,rbase
				332		:	func_rom_io_display_test	=	32'h001002c4;		//[530]add      r22,4
				333		:	func_rom_io_display_test	=	32'h204002f4;		//[534]move     r23,r20
				334		:	func_rom_io_display_test	=	32'h0ec00b62;		//[538]lil      r27,66
				335		:	func_rom_io_display_test	=	32'h0ec00347;		//[53C]lil      r26,7
				336		:	func_rom_io_display_test	=	32'h0ec00801;		//[540]lil      r0,65
				337		:	func_rom_io_display_test	=	32'h10600019;		//[544]st8      r0,r25
				338		:	func_rom_io_display_test	=	32'h10a002f3;		//[548]st32     r23,r19
				339		:	func_rom_io_display_test	=	32'h10600372;		//[54C]st8      r27,r18
				340		:	func_rom_io_display_test	=	32'h2040003e;		//[550]move     r1,rbase
				341		:	func_rom_io_display_test	=	32'h00100028;		//[554]add      r1,8
				342		:	func_rom_io_display_test	=	32'h0ee00040;		//[558]lih      r2,0x0
				343		:	func_rom_io_display_test	=	32'h0d417850;		//[55C]wl16     r2,0xbd0
				344		:	func_rom_io_display_test	=	32'h0ee003a0;		//[560]lih      rtmp,0x0
				345		:	func_rom_io_display_test	=	32'h0d416bb0;		//[564]wl16     rtmp,0xb50
				346		:	func_rom_io_display_test	=	32'h207003e2;		//[568]movepc   rret,8
				347		:	func_rom_io_display_test	=	32'h144003a0;		//[56C]b        rtmp,#al
				348		:	func_rom_io_display_test	=	32'h10a002fe;		//[570]st32     r23,rbase
				349		:	func_rom_io_display_test	=	32'h2040003e;		//[574]move     r1,rbase
				350		:	func_rom_io_display_test	=	32'h00100428;		//[578]add      r1,40
				351		:	func_rom_io_display_test	=	32'h2040005e;		//[57C]move     r2,rbase
				352		:	func_rom_io_display_test	=	32'h00100048;		//[580]add      r2,8
				353		:	func_rom_io_display_test	=	32'h0ee003a0;		//[584]lih      rtmp,0x0
				354		:	func_rom_io_display_test	=	32'h0d4143b0;		//[588]wl16     rtmp,0xa10
				355		:	func_rom_io_display_test	=	32'h207003e2;		//[58C]movepc   rret,8
				356		:	func_rom_io_display_test	=	32'h144003a0;		//[590]b        rtmp,#al
				357		:	func_rom_io_display_test	=	32'h0ee00260;		//[594]lih      r19,0x0
				358		:	func_rom_io_display_test	=	32'h0d4e8a68;		//[598]wl16     r19,0x7448
				359		:	func_rom_io_display_test	=	32'h20400053;		//[59C]move     r2,r19
				360		:	func_rom_io_display_test	=	32'h0ec00021;		//[5A0]lil      r1,1
				361		:	func_rom_io_display_test	=	32'h00d00000;		//[5A4]cmp      r0,0
				362		:	func_rom_io_display_test	=	32'h14310002;		//[5A8]br       5b0 <start+0x1d0>,#eq
				363		:	func_rom_io_display_test	=	32'h0ec00020;		//[5AC]lil      r1,0
				364		:	func_rom_io_display_test	=	32'h10a00022;		//[5B0]st32     r1,r2
				365		:	func_rom_io_display_test	=	32'h10a00356;		//[5B4]st32     r26,r22
				366		:	func_rom_io_display_test	=	32'h0ec00022;		//[5B8]lil      r1,2
				367		:	func_rom_io_display_test	=	32'h0ec00043;		//[5BC]lil      r2,3
				368		:	func_rom_io_display_test	=	32'h20400076;		//[5C0]move     r3,r22
				369		:	func_rom_io_display_test	=	32'h0ee003a0;		//[5C4]lih      rtmp,0x0
				370		:	func_rom_io_display_test	=	32'h0d411fb0;		//[5C8]wl16     rtmp,0x8f0
				371		:	func_rom_io_display_test	=	32'h207003e2;		//[5CC]movepc   rret,8
				372		:	func_rom_io_display_test	=	32'h144003a0;		//[5D0]b        rtmp,#al
				373		:	func_rom_io_display_test	=	32'h0ee00020;		//[5D4]lih      r1,0x0
				374		:	func_rom_io_display_test	=	32'h0d4e7020;		//[5D8]wl16     r1,0x7380
				375		:	func_rom_io_display_test	=	32'h0ee00040;		//[5DC]lih      r2,0x0
				376		:	func_rom_io_display_test	=	32'h0d498850;		//[5E0]wl16     r2,0x4c50
				377		:	func_rom_io_display_test	=	32'h0ec00063;		//[5E4]lil      r3,3
				378		:	func_rom_io_display_test	=	32'h10400096;		//[5E8]ld32     r4,r22
				379		:	func_rom_io_display_test	=	32'h0ee003a0;		//[5EC]lih      rtmp,0x0
				380		:	func_rom_io_display_test	=	32'h0d4123b0;		//[5F0]wl16     rtmp,0x910
				381		:	func_rom_io_display_test	=	32'h207003e2;		//[5F4]movepc   rret,8
				382		:	func_rom_io_display_test	=	32'h144003a0;		//[5F8]b        rtmp,#al
				383		:	func_rom_io_display_test	=	32'h10400038;		//[5FC]ld32     r1,r24
				384		:	func_rom_io_display_test	=	32'h0ee003a0;		//[600]lih      rtmp,0x0
				385		:	func_rom_io_display_test	=	32'h0d4023b0;		//[604]wl16     rtmp,0x110
				386		:	func_rom_io_display_test	=	32'h207003e2;		//[608]movepc   rret,8
				387		:	func_rom_io_display_test	=	32'h144003a0;		//[60C]b        rtmp,#al
				388		:	func_rom_io_display_test	=	32'h10000032;		//[610]ld8      r1,r18
				389		:	func_rom_io_display_test	=	32'h03800001;		//[614]sext8    r0,r1
				390		:	func_rom_io_display_test	=	32'h00d00800;		//[618]cmp      r0,64
				391		:	func_rom_io_display_test	=	32'h143f002c;		//[61C]br       6cc <start+0x2ec>,#seu
				392		:	func_rom_io_display_test	=	32'h0ec00a01;		//[620]lil      r16,65
				393		:	func_rom_io_display_test	=	32'h20400230;		//[624]move     r17,r16
				394		:	func_rom_io_display_test	=	32'h0ee002a0;		//[628]lih      r21,0x0
				395		:	func_rom_io_display_test	=	32'h0d4e6ea8;		//[62C]wl16     r21,0x7368
				396		:	func_rom_io_display_test	=	32'h14300008;		//[630]br       650 <start+0x270>,#al
				397		:	func_rom_io_display_test	=	32'h00100221;		//[634]add      r17,1
				398		:	func_rom_io_display_test	=	32'h03800231;		//[638]sext8    r17,r17
				399		:	func_rom_io_display_test	=	32'h00100201;		//[63C]add      r16,1
				400		:	func_rom_io_display_test	=	32'h10000052;		//[640]ld8      r2,r18
				401		:	func_rom_io_display_test	=	32'h03800002;		//[644]sext8    r0,r2
				402		:	func_rom_io_display_test	=	32'h00c00011;		//[648]cmp      r0,r17
				403		:	func_rom_io_display_test	=	32'h143d0020;		//[64C]br       6cc <start+0x2ec>,#su
				404		:	func_rom_io_display_test	=	32'h20400030;		//[650]move     r1,r16
				405		:	func_rom_io_display_test	=	32'h0ec00843;		//[654]lil      r2,67
				406		:	func_rom_io_display_test	=	32'h0ee003a0;		//[658]lih      rtmp,0x0
				407		:	func_rom_io_display_test	=	32'h0d413bb0;		//[65C]wl16     rtmp,0x9d0
				408		:	func_rom_io_display_test	=	32'h207003e2;		//[660]movepc   rret,8
				409		:	func_rom_io_display_test	=	32'h144003a0;		//[664]b        rtmp,#al
				410		:	func_rom_io_display_test	=	32'h1040003e;		//[668]ld32     r1,rbase
				411		:	func_rom_io_display_test	=	32'h00c00001;		//[66C]cmp      r0,r1
				412		:	func_rom_io_display_test	=	32'h1432fff1;		//[670]br       634 <start+0x254>,#neq
				413		:	func_rom_io_display_test	=	32'h0ec00020;		//[674]lil      r1,0
				414		:	func_rom_io_display_test	=	32'h2040005e;		//[678]move     r2,rbase
				415		:	func_rom_io_display_test	=	32'h0ee003a0;		//[67C]lih      rtmp,0x0
				416		:	func_rom_io_display_test	=	32'h0d410fa0;		//[680]wl16     rtmp,0x860
				417		:	func_rom_io_display_test	=	32'h207003e2;		//[684]movepc   rret,8
				418		:	func_rom_io_display_test	=	32'h144003a0;		//[688]b        rtmp,#al
				419		:	func_rom_io_display_test	=	32'h2040003e;		//[68C]move     r1,rbase
				420		:	func_rom_io_display_test	=	32'h00100028;		//[690]add      r1,8
				421		:	func_rom_io_display_test	=	32'h0ee00040;		//[694]lih      r2,0x0
				422		:	func_rom_io_display_test	=	32'h0d417c50;		//[698]wl16     r2,0xbf0
				423		:	func_rom_io_display_test	=	32'h0ee003a0;		//[69C]lih      rtmp,0x0
				424		:	func_rom_io_display_test	=	32'h0d416bb0;		//[6A0]wl16     rtmp,0xb50
				425		:	func_rom_io_display_test	=	32'h207003e2;		//[6A4]movepc   rret,8
				426		:	func_rom_io_display_test	=	32'h144003a0;		//[6A8]b        rtmp,#al
				427		:	func_rom_io_display_test	=	32'h10a00295;		//[6AC]st32     r20,r21
				428		:	func_rom_io_display_test	=	32'h00100221;		//[6B0]add      r17,1
				429		:	func_rom_io_display_test	=	32'h03800231;		//[6B4]sext8    r17,r17
				430		:	func_rom_io_display_test	=	32'h00100201;		//[6B8]add      r16,1
				431		:	func_rom_io_display_test	=	32'h10000052;		//[6BC]ld8      r2,r18
				432		:	func_rom_io_display_test	=	32'h03800002;		//[6C0]sext8    r0,r2
				433		:	func_rom_io_display_test	=	32'h00c00011;		//[6C4]cmp      r0,r17
				434		:	func_rom_io_display_test	=	32'h143cffe2;		//[6C8]br       650 <start+0x270>,#seo
				435		:	func_rom_io_display_test	=	32'h00100281;		//[6CC]add      r20,1
				436		:	func_rom_io_display_test	=	32'h00d00e85;		//[6D0]cmp      r20,101
				437		:	func_rom_io_display_test	=	32'h1432ff9b;		//[6D4]br       540 <start+0x160>,#neq
				438		:	func_rom_io_display_test	=	32'h0ee003a0;		//[6D8]lih      rtmp,0x0
				439		:	func_rom_io_display_test	=	32'h0d415bb0;		//[6DC]wl16     rtmp,0xad0
				440		:	func_rom_io_display_test	=	32'h207003e2;		//[6E0]movepc   rret,8
				441		:	func_rom_io_display_test	=	32'h144003a0;		//[6E4]b        rtmp,#al
				442		:	func_rom_io_display_test	=	32'h0ee00020;		//[6E8]lih      r1,0x0
				443		:	func_rom_io_display_test	=	32'h0d4e6c20;		//[6EC]wl16     r1,0x7360
				444		:	func_rom_io_display_test	=	32'h10a00001;		//[6F0]st32     r0,r1
				445		:	func_rom_io_display_test	=	32'h0ec00828;		//[6F4]lil      r1,72
				446		:	func_rom_io_display_test	=	32'h0000003e;		//[6F8]add      r1,rbase
				447		:	func_rom_io_display_test	=	32'h10400021;		//[6FC]ld32     r1,r1
				448		:	func_rom_io_display_test	=	32'h10400061;		//[700]ld32     r3,r1
				449		:	func_rom_io_display_test	=	32'h0ee00020;		//[704]lih      r1,0x0
				450		:	func_rom_io_display_test	=	32'h0d498820;		//[708]wl16     r1,0x4c40
				451		:	func_rom_io_display_test	=	32'h20400040;		//[70C]move     r2,r0
				452		:	func_rom_io_display_test	=	32'h00200043;		//[710]sub      r2,r3
				453		:	func_rom_io_display_test	=	32'h10a00041;		//[714]st32     r2,r1
				454		:	func_rom_io_display_test	=	32'h0ee02020;		//[718]lih      r1,0x100
				455		:	func_rom_io_display_test	=	32'h10a00061;		//[71C]st32     r3,r1
				456		:	func_rom_io_display_test	=	32'h0ee02020;		//[720]lih      r1,0x100
				457		:	func_rom_io_display_test	=	32'h0d400024;		//[724]wl16     r1,0x4
				458		:	func_rom_io_display_test	=	32'h10a00001;		//[728]st32     r0,r1
				459		:	func_rom_io_display_test	=	32'h0ee02000;		//[72C]lih      r0,0x100
				460		:	func_rom_io_display_test	=	32'h0d400008;		//[730]wl16     r0,0x8
				461		:	func_rom_io_display_test	=	32'h10a00040;		//[734]st32     r2,r0
				462		:	func_rom_io_display_test	=	32'h0ee02000;		//[738]lih      r0,0x100
				463		:	func_rom_io_display_test	=	32'h0d40000c;		//[73C]wl16     r0,0xc
				464		:	func_rom_io_display_test	=	32'h0ec00c24;		//[740]lil      r1,100
				465		:	func_rom_io_display_test	=	32'h10a00020;		//[744]st32     r1,r0
				466		:	func_rom_io_display_test	=	32'h180003a0;		//[748]srspr    rtmp
				467		:	func_rom_io_display_test	=	32'h00100bac;		//[74C]add      rtmp,76
				468		:	func_rom_io_display_test	=	32'h1c0003a0;		//[750]srspw    rtmp
				469		:	func_rom_io_display_test	=	32'h120003e0;		//[754]pop      rret
				470		:	func_rom_io_display_test	=	32'h12000360;		//[758]pop      r27
				471		:	func_rom_io_display_test	=	32'h12000340;		//[75C]pop      r26
				472		:	func_rom_io_display_test	=	32'h12000320;		//[760]pop      r25
				473		:	func_rom_io_display_test	=	32'h12000300;		//[764]pop      r24
				474		:	func_rom_io_display_test	=	32'h120002e0;		//[768]pop      r23
				475		:	func_rom_io_display_test	=	32'h120002c0;		//[76C]pop      r22
				476		:	func_rom_io_display_test	=	32'h120002a0;		//[770]pop      r21
				477		:	func_rom_io_display_test	=	32'h12000280;		//[774]pop      r20
				478		:	func_rom_io_display_test	=	32'h12000260;		//[778]pop      r19
				479		:	func_rom_io_display_test	=	32'h12000240;		//[77C]pop      r18
				480		:	func_rom_io_display_test	=	32'h12000220;		//[780]pop      r17
				481		:	func_rom_io_display_test	=	32'h12000200;		//[784]pop      r16
				482		:	func_rom_io_display_test	=	32'h120003c0;		//[788]pop      rbase
				483		:	func_rom_io_display_test	=	32'h144003e0;		//[78C]b        rret,#al
				484		:	func_rom_io_display_test	=	32'h110003c0;		//[790]push     rbase
				485		:	func_rom_io_display_test	=	32'h180003c0;		//[794]srspr    rbase
				486		:	func_rom_io_display_test	=	32'h0ee00020;		//[798]lih      r1,0x0
				487		:	func_rom_io_display_test	=	32'h0d4e8828;		//[79C]wl16     r1,0x7448
				488		:	func_rom_io_display_test	=	32'h0ee00000;		//[7A0]lih      r0,0x0
				489		:	func_rom_io_display_test	=	32'h0d4e6c0c;		//[7A4]wl16     r0,0x736c
				490		:	func_rom_io_display_test	=	32'h10000000;		//[7A8]ld8      r0,r0
				491		:	func_rom_io_display_test	=	32'h0ec00841;		//[7AC]lil      r2,65
				492		:	func_rom_io_display_test	=	32'h0c400002;		//[7B0]xor      r0,r2
				493		:	func_rom_io_display_test	=	32'h0e700000;		//[7B4]get8     r0,0x0
				494		:	func_rom_io_display_test	=	32'h0010fc1f;		//[7B8]add      r0,-1
				495		:	func_rom_io_display_test	=	32'h0830001f;		//[7BC]shr      r0,0x1f
				496		:	func_rom_io_display_test	=	32'h10400041;		//[7C0]ld32     r2,r1
				497		:	func_rom_io_display_test	=	32'h0c200002;		//[7C4]or       r0,r2
				498		:	func_rom_io_display_test	=	32'h10a00001;		//[7C8]st32     r0,r1
				499		:	func_rom_io_display_test	=	32'h0ee00000;		//[7CC]lih      r0,0x0
				500		:	func_rom_io_display_test	=	32'h0d4e6c0d;		//[7D0]wl16     r0,0x736d
				501		:	func_rom_io_display_test	=	32'h0ec00822;		//[7D4]lil      r1,66
				502		:	func_rom_io_display_test	=	32'h10600020;		//[7D8]st8      r1,r0
				503		:	func_rom_io_display_test	=	32'h120003c0;		//[7DC]pop      rbase
				504		:	func_rom_io_display_test	=	32'h144003e0;		//[7E0]b        rret,#al
				508		:	func_rom_io_display_test	=	32'h110003c0;		//[7F0]push     rbase
				509		:	func_rom_io_display_test	=	32'h180003c0;		//[7F4]srspr    rbase
				510		:	func_rom_io_display_test	=	32'h0ee00000;		//[7F8]lih      r0,0x0
				511		:	func_rom_io_display_test	=	32'h0d4e6c0c;		//[7FC]wl16     r0,0x736c
				512		:	func_rom_io_display_test	=	32'h0ec00821;		//[800]lil      r1,65
				513		:	func_rom_io_display_test	=	32'h10600020;		//[804]st8      r1,r0
				514		:	func_rom_io_display_test	=	32'h0ee00000;		//[808]lih      r0,0x0
				515		:	func_rom_io_display_test	=	32'h0d4e8808;		//[80C]wl16     r0,0x7448
				516		:	func_rom_io_display_test	=	32'h0ec00020;		//[810]lil      r1,0
				517		:	func_rom_io_display_test	=	32'h10a00020;		//[814]st32     r1,r0
				518		:	func_rom_io_display_test	=	32'h120003c0;		//[818]pop      rbase
				519		:	func_rom_io_display_test	=	32'h144003e0;		//[81C]b        rret,#al
				520		:	func_rom_io_display_test	=	32'h110003c0;		//[820]push     rbase
				521		:	func_rom_io_display_test	=	32'h180003c0;		//[824]srspr    rbase
				522		:	func_rom_io_display_test	=	32'h00d00060;		//[828]cmp      r3,0
				523		:	func_rom_io_display_test	=	32'h14310009;		//[82C]br       850 <memcpy+0x30>,#eq
				524		:	func_rom_io_display_test	=	32'h00000061;		//[830]add      r3,r1
				525		:	func_rom_io_display_test	=	32'h10000082;		//[834]ld8      r4,r2
				526		:	func_rom_io_display_test	=	32'h03800004;		//[838]sext8    r0,r4
				527		:	func_rom_io_display_test	=	32'h10600001;		//[83C]st8      r0,r1
				528		:	func_rom_io_display_test	=	32'h00100021;		//[840]add      r1,1
				529		:	func_rom_io_display_test	=	32'h00100041;		//[844]add      r2,1
				530		:	func_rom_io_display_test	=	32'h00c00023;		//[848]cmp      r1,r3
				531		:	func_rom_io_display_test	=	32'h1432fffa;		//[84C]br       834 <memcpy+0x14>,#neq
				532		:	func_rom_io_display_test	=	32'h120003c0;		//[850]pop      rbase
				533		:	func_rom_io_display_test	=	32'h144003e0;		//[854]b        rret,#al
				536		:	func_rom_io_display_test	=	32'h110003c0;		//[860]push     rbase
				537		:	func_rom_io_display_test	=	32'h180003c0;		//[864]srspr    rbase
				538		:	func_rom_io_display_test	=	32'h10a00022;		//[868]st32     r1,r2
				539		:	func_rom_io_display_test	=	32'h00d00022;		//[86C]cmp      r1,2
				540		:	func_rom_io_display_test	=	32'h14310013;		//[870]br       8bc <Proc_6+0x5c>,#eq
				541		:	func_rom_io_display_test	=	32'h0ec00003;		//[874]lil      r0,3
				542		:	func_rom_io_display_test	=	32'h10a00002;		//[878]st32     r0,r2
				543		:	func_rom_io_display_test	=	32'h00d00021;		//[87C]cmp      r1,1
				544		:	func_rom_io_display_test	=	32'h14310013;		//[880]br       8cc <Proc_6+0x6c>,#eq
				545		:	func_rom_io_display_test	=	32'h00d00021;		//[884]cmp      r1,1
				546		:	func_rom_io_display_test	=	32'h14380005;		//[888]br       89c <Proc_6+0x3c>,#ueo
				547		:	func_rom_io_display_test	=	32'h0ec00000;		//[88C]lil      r0,0
				548		:	func_rom_io_display_test	=	32'h10a00002;		//[890]st32     r0,r2
				549		:	func_rom_io_display_test	=	32'h120003c0;		//[894]pop      rbase
				550		:	func_rom_io_display_test	=	32'h144003e0;		//[898]b        rret,#al
				551		:	func_rom_io_display_test	=	32'h00d00022;		//[89C]cmp      r1,2
				552		:	func_rom_io_display_test	=	32'h14310007;		//[8A0]br       8bc <Proc_6+0x5c>,#eq
				553		:	func_rom_io_display_test	=	32'h00d00024;		//[8A4]cmp      r1,4
				554		:	func_rom_io_display_test	=	32'h1432fffb;		//[8A8]br       894 <Proc_6+0x34>,#neq
				555		:	func_rom_io_display_test	=	32'h0ec00002;		//[8AC]lil      r0,2
				556		:	func_rom_io_display_test	=	32'h10a00002;		//[8B0]st32     r0,r2
				557		:	func_rom_io_display_test	=	32'h120003c0;		//[8B4]pop      rbase
				558		:	func_rom_io_display_test	=	32'h144003e0;		//[8B8]b        rret,#al
				559		:	func_rom_io_display_test	=	32'h0ec00001;		//[8BC]lil      r0,1
				560		:	func_rom_io_display_test	=	32'h10a00002;		//[8C0]st32     r0,r2
				561		:	func_rom_io_display_test	=	32'h120003c0;		//[8C4]pop      rbase
				562		:	func_rom_io_display_test	=	32'h144003e0;		//[8C8]b        rret,#al
				563		:	func_rom_io_display_test	=	32'h0ee00000;		//[8CC]lih      r0,0x0
				564		:	func_rom_io_display_test	=	32'h0d4e6c08;		//[8D0]wl16     r0,0x7368
				565		:	func_rom_io_display_test	=	32'h10400000;		//[8D4]ld32     r0,r0
				566		:	func_rom_io_display_test	=	32'h00d00c04;		//[8D8]cmp      r0,100
				567		:	func_rom_io_display_test	=	32'h143effec;		//[8DC]br       88c <Proc_6+0x2c>,#so
				568		:	func_rom_io_display_test	=	32'h120003c0;		//[8E0]pop      rbase
				569		:	func_rom_io_display_test	=	32'h144003e0;		//[8E4]b        rret,#al
				572		:	func_rom_io_display_test	=	32'h110003c0;		//[8F0]push     rbase
				573		:	func_rom_io_display_test	=	32'h180003c0;		//[8F4]srspr    rbase
				574		:	func_rom_io_display_test	=	32'h00100022;		//[8F8]add      r1,2
				575		:	func_rom_io_display_test	=	32'h00000022;		//[8FC]add      r1,r2
				576		:	func_rom_io_display_test	=	32'h10a00023;		//[900]st32     r1,r3
				577		:	func_rom_io_display_test	=	32'h120003c0;		//[904]pop      rbase
				578		:	func_rom_io_display_test	=	32'h144003e0;		//[908]b        rret,#al
				579		:	func_rom_io_display_test	=	32'h00000000;		//[90C]add      r0,r0
				580		:	func_rom_io_display_test	=	32'h110003c0;		//[910]push     rbase
				581		:	func_rom_io_display_test	=	32'h180003c0;		//[914]srspr    rbase
				582		:	func_rom_io_display_test	=	32'h204000a3;		//[918]move     r5,r3
				583		:	func_rom_io_display_test	=	32'h001000a5;		//[91C]add      r5,5
				584		:	func_rom_io_display_test	=	32'h204000e5;		//[920]move     r7,r5
				585		:	func_rom_io_display_test	=	32'h081000e2;		//[924]shl      r7,0x2
				586		:	func_rom_io_display_test	=	32'h20400101;		//[928]move     r8,r1
				587		:	func_rom_io_display_test	=	32'h00000107;		//[92C]add      r8,r7
				588		:	func_rom_io_display_test	=	32'h10a00088;		//[930]st32     r4,r8
				589		:	func_rom_io_display_test	=	32'h204000c3;		//[934]move     r6,r3
				590		:	func_rom_io_display_test	=	32'h001000c6;		//[938]add      r6,6
				591		:	func_rom_io_display_test	=	32'h081000c2;		//[93C]shl      r6,0x2
				592		:	func_rom_io_display_test	=	32'h20400001;		//[940]move     r0,r1
				593		:	func_rom_io_display_test	=	32'h00000006;		//[944]add      r0,r6
				594		:	func_rom_io_display_test	=	32'h10a00080;		//[948]st32     r4,r0
				595		:	func_rom_io_display_test	=	32'h20400003;		//[94C]move     r0,r3
				596		:	func_rom_io_display_test	=	32'h00100403;		//[950]add      r0,35
				597		:	func_rom_io_display_test	=	32'h08100002;		//[954]shl      r0,0x2
				598		:	func_rom_io_display_test	=	32'h00000001;		//[958]add      r0,r1
				599		:	func_rom_io_display_test	=	32'h10a000a0;		//[95C]st32     r5,r0
				600		:	func_rom_io_display_test	=	32'h0ec01808;		//[960]lil      r0,200
				601		:	func_rom_io_display_test	=	32'h00400005;		//[964]mull     r0,r5
				602		:	func_rom_io_display_test	=	32'h00000002;		//[968]add      r0,r2
				603		:	func_rom_io_display_test	=	32'h20400020;		//[96C]move     r1,r0
				604		:	func_rom_io_display_test	=	32'h00000027;		//[970]add      r1,r7
				605		:	func_rom_io_display_test	=	32'h10a000a1;		//[974]st32     r5,r1
				606		:	func_rom_io_display_test	=	32'h000000c0;		//[978]add      r6,r0
				607		:	func_rom_io_display_test	=	32'h10a000a6;		//[97C]st32     r5,r6
				608		:	func_rom_io_display_test	=	32'h00100064;		//[980]add      r3,4
				609		:	func_rom_io_display_test	=	32'h08100062;		//[984]shl      r3,0x2
				610		:	func_rom_io_display_test	=	32'h00000060;		//[988]add      r3,r0
				611		:	func_rom_io_display_test	=	32'h10400023;		//[98C]ld32     r1,r3
				612		:	func_rom_io_display_test	=	32'h00100021;		//[990]add      r1,1
				613		:	func_rom_io_display_test	=	32'h10a00023;		//[994]st32     r1,r3
				614		:	func_rom_io_display_test	=	32'h10400108;		//[998]ld32     r8,r8
				615		:	func_rom_io_display_test	=	32'h0ec1f420;		//[99C]lil      r1,4000
				616		:	func_rom_io_display_test	=	32'h00000001;		//[9A0]add      r0,r1
				617		:	func_rom_io_display_test	=	32'h00000007;		//[9A4]add      r0,r7
				618		:	func_rom_io_display_test	=	32'h10a00100;		//[9A8]st32     r8,r0
				619		:	func_rom_io_display_test	=	32'h0ee00000;		//[9AC]lih      r0,0x0
				620		:	func_rom_io_display_test	=	32'h0d4e6c08;		//[9B0]wl16     r0,0x7368
				621		:	func_rom_io_display_test	=	32'h0ec00025;		//[9B4]lil      r1,5
				622		:	func_rom_io_display_test	=	32'h10a00020;		//[9B8]st32     r1,r0
				623		:	func_rom_io_display_test	=	32'h120003c0;		//[9BC]pop      rbase
				624		:	func_rom_io_display_test	=	32'h144003e0;		//[9C0]b        rret,#al
				628		:	func_rom_io_display_test	=	32'h110003c0;		//[9D0]push     rbase
				629		:	func_rom_io_display_test	=	32'h180003c0;		//[9D4]srspr    rbase
				630		:	func_rom_io_display_test	=	32'h03800001;		//[9D8]sext8    r0,r1
				631		:	func_rom_io_display_test	=	32'h03800042;		//[9DC]sext8    r2,r2
				632		:	func_rom_io_display_test	=	32'h00c00002;		//[9E0]cmp      r0,r2
				633		:	func_rom_io_display_test	=	32'h14310004;		//[9E4]br       9f4 <Func_1+0x24>,#eq
				634		:	func_rom_io_display_test	=	32'h0ec00000;		//[9E8]lil      r0,0
				635		:	func_rom_io_display_test	=	32'h120003c0;		//[9EC]pop      rbase
				636		:	func_rom_io_display_test	=	32'h144003e0;		//[9F0]b        rret,#al
				637		:	func_rom_io_display_test	=	32'h0ee00000;		//[9F4]lih      r0,0x0
				638		:	func_rom_io_display_test	=	32'h0d4e6c0c;		//[9F8]wl16     r0,0x736c
				639		:	func_rom_io_display_test	=	32'h10600020;		//[9FC]st8      r1,r0
				640		:	func_rom_io_display_test	=	32'h0ec00001;		//[A00]lil      r0,1
				641		:	func_rom_io_display_test	=	32'h120003c0;		//[A04]pop      rbase
				642		:	func_rom_io_display_test	=	32'h144003e0;		//[A08]b        rret,#al
				643		:	func_rom_io_display_test	=	32'h00000000;		//[A0C]add      r0,r0
				644		:	func_rom_io_display_test	=	32'h110003c0;		//[A10]push     rbase
				645		:	func_rom_io_display_test	=	32'h110003e0;		//[A14]push     rret
				646		:	func_rom_io_display_test	=	32'h180003c0;		//[A18]srspr    rbase
				647		:	func_rom_io_display_test	=	32'h0ee00000;		//[A1C]lih      r0,0x0
				648		:	func_rom_io_display_test	=	32'h0d4e6c0c;		//[A20]wl16     r0,0x736c
				649		:	func_rom_io_display_test	=	32'h10000080;		//[A24]ld8      r4,r0
				650		:	func_rom_io_display_test	=	32'h03800064;		//[A28]sext8    r3,r4
				651		:	func_rom_io_display_test	=	32'h204000a2;		//[A2C]move     r5,r2
				652		:	func_rom_io_display_test	=	32'h001000a3;		//[A30]add      r5,3
				653		:	func_rom_io_display_test	=	32'h20400081;		//[A34]move     r4,r1
				654		:	func_rom_io_display_test	=	32'h00100082;		//[A38]add      r4,2
				655		:	func_rom_io_display_test	=	32'h100000a5;		//[A3C]ld8      r5,r5
				656		:	func_rom_io_display_test	=	32'h038000a5;		//[A40]sext8    r5,r5
				657		:	func_rom_io_display_test	=	32'h10000084;		//[A44]ld8      r4,r4
				658		:	func_rom_io_display_test	=	32'h03800084;		//[A48]sext8    r4,r4
				659		:	func_rom_io_display_test	=	32'h00c000a4;		//[A4C]cmp      r5,r4
				660		:	func_rom_io_display_test	=	32'h14310014;		//[A50]br       aa0 <Func_2+0x90>,#eq
				661		:	func_rom_io_display_test	=	32'h10600060;		//[A54]st8      r3,r0
				662		:	func_rom_io_display_test	=	32'h0ee003a0;		//[A58]lih      rtmp,0x0
				663		:	func_rom_io_display_test	=	32'h0d4163a0;		//[A5C]wl16     rtmp,0xb00
				664		:	func_rom_io_display_test	=	32'h207003e2;		//[A60]movepc   rret,8
				665		:	func_rom_io_display_test	=	32'h144003a0;		//[A64]b        rtmp,#al
				666		:	func_rom_io_display_test	=	32'h00d00000;		//[A68]cmp      r0,0
				667		:	func_rom_io_display_test	=	32'h143f0009;		//[A6C]br       a90 <Func_2+0x80>,#seu
				668		:	func_rom_io_display_test	=	32'h0ee00000;		//[A70]lih      r0,0x0
				669		:	func_rom_io_display_test	=	32'h0d4e6c08;		//[A74]wl16     r0,0x7368
				670		:	func_rom_io_display_test	=	32'h0ec0002a;		//[A78]lil      r1,10
				671		:	func_rom_io_display_test	=	32'h10a00020;		//[A7C]st32     r1,r0
				672		:	func_rom_io_display_test	=	32'h0ec00001;		//[A80]lil      r0,1
				673		:	func_rom_io_display_test	=	32'h120003e0;		//[A84]pop      rret
				674		:	func_rom_io_display_test	=	32'h120003c0;		//[A88]pop      rbase
				675		:	func_rom_io_display_test	=	32'h144003e0;		//[A8C]b        rret,#al
				676		:	func_rom_io_display_test	=	32'h0ec00000;		//[A90]lil      r0,0
				677		:	func_rom_io_display_test	=	32'h120003e0;		//[A94]pop      rret
				678		:	func_rom_io_display_test	=	32'h120003c0;		//[A98]pop      rbase
				679		:	func_rom_io_display_test	=	32'h144003e0;		//[A9C]b        rret,#al
				680		:	func_rom_io_display_test	=	32'h14300000;		//[AA0]br       aa0 <Func_2+0x90>,#al
				684		:	func_rom_io_display_test	=	32'h110003c0;		//[AB0]push     rbase
				685		:	func_rom_io_display_test	=	32'h180003c0;		//[AB4]srspr    rbase
				686		:	func_rom_io_display_test	=	32'h0ec00001;		//[AB8]lil      r0,1
				687		:	func_rom_io_display_test	=	32'h00d00022;		//[ABC]cmp      r1,2
				688		:	func_rom_io_display_test	=	32'h14310002;		//[AC0]br       ac8 <Func_3+0x18>,#eq
				689		:	func_rom_io_display_test	=	32'h0ec00000;		//[AC4]lil      r0,0
				690		:	func_rom_io_display_test	=	32'h120003c0;		//[AC8]pop      rbase
				691		:	func_rom_io_display_test	=	32'h144003e0;		//[ACC]b        rret,#al
				692		:	func_rom_io_display_test	=	32'h110003c0;		//[AD0]push     rbase
				693		:	func_rom_io_display_test	=	32'h180003c0;		//[AD4]srspr    rbase
				694		:	func_rom_io_display_test	=	32'h1a800000;		//[AD8]srfrcr
				695		:	func_rom_io_display_test	=	32'h1ac00000;		//[ADC]srfrchr  r0
				696		:	func_rom_io_display_test	=	32'h1aa00020;		//[AE0]srfrclr  r1
				697		:	func_rom_io_display_test	=	32'h08300030;		//[AE4]shr      r1,0x10
				698		:	func_rom_io_display_test	=	32'h08100010;		//[AE8]shl      r0,0x10
				699		:	func_rom_io_display_test	=	32'h0c200001;		//[AEC]or       r0,r1
				700		:	func_rom_io_display_test	=	32'h120003c0;		//[AF0]pop      rbase
				701		:	func_rom_io_display_test	=	32'h144003e0;		//[AF4]b        rret,#al
				704		:	func_rom_io_display_test	=	32'h110003c0;		//[B00]push     rbase
				705		:	func_rom_io_display_test	=	32'h180003c0;		//[B04]srspr    rbase
				706		:	func_rom_io_display_test	=	32'h10000001;		//[B08]ld8      r0,r1
				707		:	func_rom_io_display_test	=	32'h00100021;		//[B0C]add      r1,1
				708		:	func_rom_io_display_test	=	32'h10000062;		//[B10]ld8      r3,r2
				709		:	func_rom_io_display_test	=	32'h00100041;		//[B14]add      r2,1
				710		:	func_rom_io_display_test	=	32'h00d00000;		//[B18]cmp      r0,0
				711		:	func_rom_io_display_test	=	32'h14310006;		//[B1C]br       b34 <strcmp+0x34>,#eq
				712		:	func_rom_io_display_test	=	32'h00c00003;		//[B20]cmp      r0,r3
				713		:	func_rom_io_display_test	=	32'h1431fff9;		//[B24]br       b08 <strcmp+0x8>,#eq
				714		:	func_rom_io_display_test	=	32'h00200003;		//[B28]sub      r0,r3
				715		:	func_rom_io_display_test	=	32'h120003c0;		//[B2C]pop      rbase
				716		:	func_rom_io_display_test	=	32'h144003e0;		//[B30]b        rret,#al
				717		:	func_rom_io_display_test	=	32'h20400003;		//[B34]move     r0,r3
				718		:	func_rom_io_display_test	=	32'h01200000;		//[B38]neg      r0
				719		:	func_rom_io_display_test	=	32'h120003c0;		//[B3C]pop      rbase
				720		:	func_rom_io_display_test	=	32'h144003e0;		//[B40]b        rret,#al
				724		:	func_rom_io_display_test	=	32'h110003c0;		//[B50]push     rbase
				725		:	func_rom_io_display_test	=	32'h180003c0;		//[B54]srspr    rbase
				726		:	func_rom_io_display_test	=	32'h20400001;		//[B58]move     r0,r1
				727		:	func_rom_io_display_test	=	32'h204000a1;		//[B5C]move     r5,r1
				728		:	func_rom_io_display_test	=	32'h002000a2;		//[B60]sub      r5,r2
				729		:	func_rom_io_display_test	=	32'h10000022;		//[B64]ld8      r1,r2
				730		:	func_rom_io_display_test	=	32'h03800061;		//[B68]sext8    r3,r1
				731		:	func_rom_io_display_test	=	32'h20400082;		//[B6C]move     r4,r2
				732		:	func_rom_io_display_test	=	32'h00000085;		//[B70]add      r4,r5
				733		:	func_rom_io_display_test	=	32'h10600064;		//[B74]st8      r3,r4
				734		:	func_rom_io_display_test	=	32'h00100041;		//[B78]add      r2,1
				735		:	func_rom_io_display_test	=	32'h00d00060;		//[B7C]cmp      r3,0
				736		:	func_rom_io_display_test	=	32'h1432fff9;		//[B80]br       b64 <strcpy+0x14>,#neq
				737		:	func_rom_io_display_test	=	32'h120003c0;		//[B84]pop      rbase
				738		:	func_rom_io_display_test	=	32'h144003e0;		//[B88]b        rret,#al
				739		:	func_rom_io_display_test	=	32'h00000000;		//[B8C]add      r0,r0
				740		:	func_rom_io_display_test	=	32'h44485259;		//[B90]*unknown*
				741		:	func_rom_io_display_test	=	32'h53544f4e;		//[B94]*unknown*
				742		:	func_rom_io_display_test	=	32'h45205052;		//[B98]*unknown*
				743		:	func_rom_io_display_test	=	32'h4f475241;		//[B9C]*unknown*
				744		:	func_rom_io_display_test	=	32'h4d2c2053;		//[BA0]*unknown*
				745		:	func_rom_io_display_test	=	32'h4f4d4520;		//[BA4]*unknown*
				746		:	func_rom_io_display_test	=	32'h53545249;		//[BA8]*unknown*
				747		:	func_rom_io_display_test	=	32'h4e470000;		//[BAC]*unknown*
				748		:	func_rom_io_display_test	=	32'h44485259;		//[BB0]*unknown*
				749		:	func_rom_io_display_test	=	32'h53544f4e;		//[BB4]*unknown*
				750		:	func_rom_io_display_test	=	32'h45205052;		//[BB8]*unknown*
				751		:	func_rom_io_display_test	=	32'h4f475241;		//[BBC]*unknown*
				752		:	func_rom_io_display_test	=	32'h4d2c2031;		//[BC0]*unknown*
				753		:	func_rom_io_display_test	=	32'h27535420;		//[BC4]*unknown*
				754		:	func_rom_io_display_test	=	32'h53545249;		//[BC8]*unknown*
				755		:	func_rom_io_display_test	=	32'h4e470000;		//[BCC]*unknown*
				756		:	func_rom_io_display_test	=	32'h44485259;		//[BD0]*unknown*
				757		:	func_rom_io_display_test	=	32'h53544f4e;		//[BD4]*unknown*
				758		:	func_rom_io_display_test	=	32'h45205052;		//[BD8]*unknown*
				759		:	func_rom_io_display_test	=	32'h4f475241;		//[BDC]*unknown*
				760		:	func_rom_io_display_test	=	32'h4d2c2032;		//[BE0]*unknown*
				761		:	func_rom_io_display_test	=	32'h274e4420;		//[BE4]*unknown*
				762		:	func_rom_io_display_test	=	32'h53545249;		//[BE8]*unknown*
				763		:	func_rom_io_display_test	=	32'h4e470000;		//[BEC]*unknown*
				764		:	func_rom_io_display_test	=	32'h44485259;		//[BF0]*unknown*
				765		:	func_rom_io_display_test	=	32'h53544f4e;		//[BF4]*unknown*
				766		:	func_rom_io_display_test	=	32'h45205052;		//[BF8]*unknown*
				767		:	func_rom_io_display_test	=	32'h4f475241;		//[BFC]*unknown*
				768		:	func_rom_io_display_test	=	32'h4d2c2033;		//[C00]*unknown*
				769		:	func_rom_io_display_test	=	32'h27524420;		//[C04]*unknown*
				770		:	func_rom_io_display_test	=	32'h53545249;		//[C08]*unknown*
				771		:	func_rom_io_display_test	=	32'h4e470000;		//[C0C]*unknown*
				4868		:	func_rom_io_display_test	=	32'h52656769;		//[4C10] *unknown*
				4869		:	func_rom_io_display_test	=	32'h73746572;		//[4C14] *unknown*
				4870		:	func_rom_io_display_test	=	32'h206f7074;		//[4C18] *unknown*
				4871		:	func_rom_io_display_test	=	32'h696f6e20;		//[4C1C] *unknown*
				4872		:	func_rom_io_display_test	=	32'h73656c65;		//[4C20] *unknown*
				4873		:	func_rom_io_display_test	=	32'h63746564;		//[4C24] *unknown*
				4874		:	func_rom_io_display_test	=	32'h2e000000;		//[4C28] *unknown*
				4875		:	func_rom_io_display_test	=	32'h00000000;		//[4C2C] add      r0,r0
				4876		:	func_rom_io_display_test	=	32'h04000000;		//[4C30] *unknown*
				4880		:	func_rom_io_display_test	=	32'h00000000;		//[4C40] add      r0,r0
				7384		:	func_rom_io_display_test	=	32'h00000000;		//[7360] add      r0,r0
				7385		:	func_rom_io_display_test	=	32'h00000000;		//[7364] add      r0,r0
				7386		:	func_rom_io_display_test	=	32'h00000000;		//[7368] add      r0,r0
				7387		:	func_rom_io_display_test	=	32'h00000000;		//[736C] add      r0,r0
				7442		:	func_rom_io_display_test	=	32'h00000000;		//[7448] add      r0,r0

				default	:	func_rom_io_display_test	=	32'h20000000;	//nop
			endcase
		end
	endfunction
	
	
	
	//Output Assign
	assign		oDEBUG_VALID				=		!b_write_end || !b_wait_end;
	assign		oDEBUG_MEMIF_REQ_VALID		=		!iDEBUG_MEMIF_REQ_LOCK;
	assign		oDEBUG_MEMIF_REQ_DQM0		=		1'b0;
	assign		oDEBUG_MEMIF_REQ_DQM1		=		1'b0;
	assign		oDEBUG_MEMIF_REQ_DQM2		=		1'b0;
	assign		oDEBUG_MEMIF_REQ_DQM3		=		1'b0;
	assign		oDEBUG_MEMIF_REQ_RW			=		1'b1;	//0:Read 1:Write
	assign		oDEBUG_MEMIF_REQ_ADDR		=		b_write_counter[24:0];
	assign		oDEBUG_MEMIF_REQ_DATA		=		func_rom_io_display_test(b_write_counter);//func_rom(b_write_counter);//func_rom_sysreg_test(b_write_counter);//
	
endmodule


`default_nettype wire
