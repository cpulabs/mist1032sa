library verilog;
use verilog.vl_types.all;
entity altparallel_flash_loader is
    generic(
        EXTRA_ADDR_BYTE : integer := 0;
        FEATURES_CFG    : integer := 1;
        PAGE_CLK_DIVISOR: integer := 1;
        BURST_MODE_SPANSION: integer := 0;
        ENHANCED_FLASH_PROGRAMMING: integer := 0;
        FLASH_ECC_CHECKBOX: integer := 0;
        FLASH_NRESET_COUNTER: integer := 1;
        PAGE_MODE       : integer := 0;
        NRB_ADDR        : integer := 65667072;
        BURST_MODE      : integer := 0;
        SAFE_MODE_REVERT_ADDR: integer := 0;
        US_UNIT_COUNTER : integer := 1;
        FIFO_SIZE       : integer := 16;
        CONF_DATA_WIDTH : integer := 1;
        CONF_WAIT_TIMER_WIDTH: integer := 14;
        NFLASH_MFC      : string  := "NUMONYX";
        OPTION_BITS_START_ADDRESS: integer := 0;
        SAFE_MODE_RETRY : integer := 1;
        DCLK_DIVISOR    : integer := 1;
        FLASH_TYPE      : string  := "CFI_FLASH";
        N_FLASH         : integer := 1;
        FLASH_BURST_EXTRA_CYCLE: integer := 0;
        TRISTATE_CHECKBOX: integer := 0;
        QFLASH_MFC      : string  := "ALTERA";
        FEATURES_PGM    : integer := 1;
        DISABLE_CRC_CHECKBOX: integer := 0;
        FLASH_DATA_WIDTH: integer := 16;
        RSU_WATCHDOG_COUNTER: integer := 100000000;
        PFL_RSU_WATCHDOG_ENABLED: integer := 0;
        SAFE_MODE_HALT  : integer := 0;
        ADDR_WIDTH      : integer := 20;
        NAND_SIZE       : integer := 67108864;
        NORMAL_MODE     : integer := 1;
        FLASH_NRESET_CHECKBOX: integer := 0;
        SAFE_MODE_REVERT: integer := 0;
        LPM_TYPE        : string  := "ALTPARALLEL_FLASH_LOADER";
        AUTO_RESTART    : string  := "OFF";
        CLK_DIVISOR     : integer := 1;
        BURST_MODE_INTEL: integer := 0;
        BURST_MODE_NUMONYX: integer := 0;
        DECOMPRESSOR_MODE: string  := "NONE";
        PFL_QUAD_IO_FLASH_IR_BITS: integer := 8;
        PFL_CFI_FLASH_IR_BITS: integer := 5;
        PFL_NAND_FLASH_IR_BITS: integer := 4;
        N_FLASH_BITS    : integer := 4
    );
    port(
        flash_nce       : out    vl_logic_vector;
        fpga_data       : out    vl_logic_vector;
        fpga_dclk       : out    vl_logic;
        fpga_nstatus    : in     vl_logic;
        flash_ale       : out    vl_logic;
        pfl_clk         : in     vl_logic;
        fpga_nconfig    : out    vl_logic;
        flash_io2       : inout  vl_logic_vector;
        flash_sck       : out    vl_logic_vector;
        flash_noe       : out    vl_logic;
        flash_nwe       : out    vl_logic;
        pfl_watchdog_error: out    vl_logic;
        pfl_reset_watchdog: in     vl_logic;
        fpga_conf_done  : in     vl_logic;
        flash_rdy       : in     vl_logic;
        pfl_flash_access_granted: in     vl_logic;
        pfl_nreconfigure: in     vl_logic;
        flash_cle       : out    vl_logic;
        flash_nreset    : out    vl_logic;
        flash_io0       : inout  vl_logic_vector;
        pfl_nreset      : in     vl_logic;
        flash_data      : inout  vl_logic_vector;
        flash_io1       : inout  vl_logic_vector;
        flash_nadv      : out    vl_logic;
        flash_clk       : out    vl_logic;
        flash_io3       : inout  vl_logic_vector;
        flash_io        : inout  vl_logic_vector(7 downto 0);
        flash_addr      : out    vl_logic_vector;
        pfl_flash_access_request: out    vl_logic;
        flash_ncs       : out    vl_logic_vector;
        fpga_pgm        : in     vl_logic_vector(2 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of EXTRA_ADDR_BYTE : constant is 1;
    attribute mti_svvh_generic_type of FEATURES_CFG : constant is 1;
    attribute mti_svvh_generic_type of PAGE_CLK_DIVISOR : constant is 1;
    attribute mti_svvh_generic_type of BURST_MODE_SPANSION : constant is 1;
    attribute mti_svvh_generic_type of ENHANCED_FLASH_PROGRAMMING : constant is 1;
    attribute mti_svvh_generic_type of FLASH_ECC_CHECKBOX : constant is 1;
    attribute mti_svvh_generic_type of FLASH_NRESET_COUNTER : constant is 1;
    attribute mti_svvh_generic_type of PAGE_MODE : constant is 1;
    attribute mti_svvh_generic_type of NRB_ADDR : constant is 1;
    attribute mti_svvh_generic_type of BURST_MODE : constant is 1;
    attribute mti_svvh_generic_type of SAFE_MODE_REVERT_ADDR : constant is 1;
    attribute mti_svvh_generic_type of US_UNIT_COUNTER : constant is 1;
    attribute mti_svvh_generic_type of FIFO_SIZE : constant is 1;
    attribute mti_svvh_generic_type of CONF_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CONF_WAIT_TIMER_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NFLASH_MFC : constant is 1;
    attribute mti_svvh_generic_type of OPTION_BITS_START_ADDRESS : constant is 1;
    attribute mti_svvh_generic_type of SAFE_MODE_RETRY : constant is 1;
    attribute mti_svvh_generic_type of DCLK_DIVISOR : constant is 1;
    attribute mti_svvh_generic_type of FLASH_TYPE : constant is 1;
    attribute mti_svvh_generic_type of N_FLASH : constant is 1;
    attribute mti_svvh_generic_type of FLASH_BURST_EXTRA_CYCLE : constant is 1;
    attribute mti_svvh_generic_type of TRISTATE_CHECKBOX : constant is 1;
    attribute mti_svvh_generic_type of QFLASH_MFC : constant is 1;
    attribute mti_svvh_generic_type of FEATURES_PGM : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_CRC_CHECKBOX : constant is 1;
    attribute mti_svvh_generic_type of FLASH_DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of RSU_WATCHDOG_COUNTER : constant is 1;
    attribute mti_svvh_generic_type of PFL_RSU_WATCHDOG_ENABLED : constant is 1;
    attribute mti_svvh_generic_type of SAFE_MODE_HALT : constant is 1;
    attribute mti_svvh_generic_type of ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NAND_SIZE : constant is 1;
    attribute mti_svvh_generic_type of NORMAL_MODE : constant is 1;
    attribute mti_svvh_generic_type of FLASH_NRESET_CHECKBOX : constant is 1;
    attribute mti_svvh_generic_type of SAFE_MODE_REVERT : constant is 1;
    attribute mti_svvh_generic_type of LPM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of AUTO_RESTART : constant is 1;
    attribute mti_svvh_generic_type of CLK_DIVISOR : constant is 1;
    attribute mti_svvh_generic_type of BURST_MODE_INTEL : constant is 1;
    attribute mti_svvh_generic_type of BURST_MODE_NUMONYX : constant is 1;
    attribute mti_svvh_generic_type of DECOMPRESSOR_MODE : constant is 1;
    attribute mti_svvh_generic_type of PFL_QUAD_IO_FLASH_IR_BITS : constant is 1;
    attribute mti_svvh_generic_type of PFL_CFI_FLASH_IR_BITS : constant is 1;
    attribute mti_svvh_generic_type of PFL_NAND_FLASH_IR_BITS : constant is 1;
    attribute mti_svvh_generic_type of N_FLASH_BITS : constant is 1;
end altparallel_flash_loader;
