library verilog;
use verilog.vl_types.all;
entity reservation_alu3_entry is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iREMOVE_VALID   : in     vl_logic;
        iREGISTER_VALID : in     vl_logic;
        iREGISTER_CMD   : in     vl_logic_vector(4 downto 0);
        iREGISTER_SYS_LDST: in     vl_logic;
        iREGISTER_LDST  : in     vl_logic;
        iREGISTER_SOURCE0_VALID: in     vl_logic;
        iREGISTER_SOURCE0_SYSREG: in     vl_logic;
        iREGISTER_SOURCE0: in     vl_logic_vector(31 downto 0);
        iREGISTER_SOURCE1_VALID: in     vl_logic;
        iREGISTER_SOURCE1_SYSREG: in     vl_logic;
        iREGISTER_SOURCE1: in     vl_logic_vector(31 downto 0);
        iREGISTER_ADV_ACTIVE: in     vl_logic;
        iREGISTER_ADV_DATA: in     vl_logic_vector(5 downto 0);
        iREGISTER_LOGIC_DEST: in     vl_logic_vector(4 downto 0);
        iREGISTER_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iREGISTER_DESTINATION_SYSREG: in     vl_logic;
        iREGISTER_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iREGISTER_PC    : in     vl_logic_vector(31 downto 0);
        iREGISTER_EX_REGIST_POINTER: in     vl_logic_vector(3 downto 0);
        iADDER_VALID    : in     vl_logic;
        iADDER_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iADDER_WRITEBACK: in     vl_logic;
        iADDER_DATA     : in     vl_logic_vector(31 downto 0);
        iMULDIV_VALID   : in     vl_logic;
        iMULDIV_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iMULDIV_WRITEBACK: in     vl_logic;
        iMULDIV_DATA    : in     vl_logic_vector(31 downto 0);
        iLDST_VALID     : in     vl_logic;
        iLDST_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iLDST_DATA      : in     vl_logic_vector(31 downto 0);
        iEX_EXECUTION_POINTER: in     vl_logic_vector(3 downto 0);
        iEXOUT_VALID    : in     vl_logic;
        oINFO_ENTRY_VALID: out    vl_logic;
        oINFO_MATCHING  : out    vl_logic;
        oINFO_CMD       : out    vl_logic_vector(4 downto 0);
        oINFO_SYS_LDST  : out    vl_logic;
        oINFO_LDST      : out    vl_logic;
        oINFO_SOURCE0_VALID: out    vl_logic;
        oINFO_SOURCE0_SYSREG: out    vl_logic;
        oINFO_SOURCE0   : out    vl_logic_vector(31 downto 0);
        oINFO_SOURCE1_VALID: out    vl_logic;
        oINFO_SOURCE1_SYSREG: out    vl_logic;
        oINFO_SOURCE1   : out    vl_logic_vector(31 downto 0);
        oINFO_ADV_ACTIVE: out    vl_logic;
        oINFO_ADV_DATA  : out    vl_logic_vector(5 downto 0);
        oINFO_LOGIC_DEST: out    vl_logic_vector(4 downto 0);
        oINFO_DESTINATION_REGNAME: out    vl_logic_vector(5 downto 0);
        oINFO_DESTINATION_SYSREG: out    vl_logic;
        oINFO_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oINFO_PC        : out    vl_logic_vector(31 downto 0)
    );
end reservation_alu3_entry;
