library verilog;
use verilog.vl_types.all;
entity scheduler2 is
    generic(
        CORE_ID         : integer := 0
    );
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iFREE_DEFAULT   : in     vl_logic;
        iFREE_RESTART   : in     vl_logic;
        iFREE_RESERVATIONSTATION: in     vl_logic;
        iFREE_SYSREG_SET_IRQ_MODE: in     vl_logic;
        iFREE_SYSREG_BACK_PREVIOUS: in     vl_logic;
        iFREE_CURRENT_PC: in     vl_logic_vector(31 downto 0);
        iFREE_REGISTER  : in     vl_logic_vector(63 downto 0);
        iCOMMIT_ENTRY_COMMIT_VECTOR: in     vl_logic_vector(63 downto 0);
        iSYSREGINFO_IOSR_VALID: in     vl_logic;
        iSYSREGINFO_IOSR: in     vl_logic_vector(31 downto 0);
        oSYSREGINFO_TIDR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_PTIDR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_PSR : out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_PPSR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_TISR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_PDTR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_IDTR: out    vl_logic_vector(31 downto 0);
        oSYSREGINFO_PPCR: out    vl_logic_vector(31 downto 0);
        iPREVIOUS_0_VALID: in     vl_logic;
        iPREVIOUS_0_SOURCE0_ACTIVE: in     vl_logic;
        iPREVIOUS_0_SOURCE1_ACTIVE: in     vl_logic;
        iPREVIOUS_0_SOURCE0_SYSREG: in     vl_logic;
        iPREVIOUS_0_SOURCE1_SYSREG: in     vl_logic;
        iPREVIOUS_0_SOURCE0_SYSREG_RENAME: in     vl_logic;
        iPREVIOUS_0_SOURCE1_SYSREG_RENAME: in     vl_logic;
        iPREVIOUS_0_ADV_ACTIVE: in     vl_logic;
        iPREVIOUS_0_DESTINATION_SYSREG: in     vl_logic;
        iPREVIOUS_0_WRITEBACK: in     vl_logic;
        iPREVIOUS_0_FLAGS_WRITEBACK: in     vl_logic;
        iPREVIOUS_0_CMD : in     vl_logic_vector(4 downto 0);
        iPREVIOUS_0_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_0_CC_AFE: in     vl_logic_vector(3 downto 0);
        iPREVIOUS_0_FLAGS_REGNAME: in     vl_logic_vector(3 downto 0);
        iPREVIOUS_0_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_0_LOGIC_DESTINATION: in     vl_logic_vector(4 downto 0);
        iPREVIOUS_0_SOURCE0: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_0_SOURCE1: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_0_ADV_DATA: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_0_SOURCE0_FLAGS: in     vl_logic;
        iPREVIOUS_0_SOURCE1_IMM: in     vl_logic;
        iPREVIOUS_0_EX_SYS_REG: in     vl_logic;
        iPREVIOUS_0_EX_SYS_LDST: in     vl_logic;
        iPREVIOUS_0_EX_LOGIC: in     vl_logic;
        iPREVIOUS_0_EX_SHIFT: in     vl_logic;
        iPREVIOUS_0_EX_ADDER: in     vl_logic;
        iPREVIOUS_0_EX_MUL: in     vl_logic;
        iPREVIOUS_0_EX_SDIV: in     vl_logic;
        iPREVIOUS_0_EX_UDIV: in     vl_logic;
        iPREVIOUS_0_EX_LDST: in     vl_logic;
        iPREVIOUS_0_EX_BRANCH: in     vl_logic;
        iPREVIOUS_1_VALID: in     vl_logic;
        iPREVIOUS_1_SOURCE0_ACTIVE: in     vl_logic;
        iPREVIOUS_1_SOURCE1_ACTIVE: in     vl_logic;
        iPREVIOUS_1_SOURCE0_SYSREG: in     vl_logic;
        iPREVIOUS_1_SOURCE1_SYSREG: in     vl_logic;
        iPREVIOUS_1_SOURCE0_SYSREG_RENAME: in     vl_logic;
        iPREVIOUS_1_SOURCE1_SYSREG_RENAME: in     vl_logic;
        iPREVIOUS_1_ADV_ACTIVE: in     vl_logic;
        iPREVIOUS_1_DESTINATION_SYSREG: in     vl_logic;
        iPREVIOUS_1_WRITEBACK: in     vl_logic;
        iPREVIOUS_1_FLAGS_WRITEBACK: in     vl_logic;
        iPREVIOUS_1_CMD : in     vl_logic_vector(4 downto 0);
        iPREVIOUS_1_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_1_CC_AFE: in     vl_logic_vector(3 downto 0);
        iPREVIOUS_1_FLAGS_REGNAME: in     vl_logic_vector(3 downto 0);
        iPREVIOUS_1_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_1_LOGIC_DESTINATION: in     vl_logic_vector(4 downto 0);
        iPREVIOUS_1_SOURCE0: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_1_SOURCE1: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_1_ADV_DATA: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_1_SOURCE0_FLAGS: in     vl_logic;
        iPREVIOUS_1_SOURCE1_IMM: in     vl_logic;
        iPREVIOUS_1_EX_SYS_REG: in     vl_logic;
        iPREVIOUS_1_EX_SYS_LDST: in     vl_logic;
        iPREVIOUS_1_EX_LOGIC: in     vl_logic;
        iPREVIOUS_1_EX_SHIFT: in     vl_logic;
        iPREVIOUS_1_EX_ADDER: in     vl_logic;
        iPREVIOUS_1_EX_MUL: in     vl_logic;
        iPREVIOUS_1_EX_SDIV: in     vl_logic;
        iPREVIOUS_1_EX_UDIV: in     vl_logic;
        iPREVIOUS_1_EX_LDST: in     vl_logic;
        iPREVIOUS_1_EX_BRANCH: in     vl_logic;
        iPREVIOUS_PC    : in     vl_logic_vector(31 downto 0);
        oPREVIOUS_LOCK  : out    vl_logic;
        oFLAG_REGISTER_0_WR: out    vl_logic;
        oFLAG_REGISTER_0_NUM: out    vl_logic_vector(3 downto 0);
        iFLAG_REGISTER_0_FULL: in     vl_logic;
        iFLAG_REGISTER_0_COUNT: in     vl_logic_vector(1 downto 0);
        oFLAG_REGISTER_1_WR: out    vl_logic;
        oFLAG_REGISTER_1_NUM: out    vl_logic_vector(3 downto 0);
        iFLAG_REGISTER_1_FULL: in     vl_logic;
        iFLAG_REGISTER_1_COUNT: in     vl_logic_vector(1 downto 0);
        oOTHER_REGISTER_0_WR: out    vl_logic;
        oOTHER_REGISTER_0_NUM: out    vl_logic_vector(5 downto 0);
        iOTHER_REGISTER_0_FULL: in     vl_logic;
        iOTHER_REGISTER_0_COUNT: in     vl_logic_vector(2 downto 0);
        oOTHER_REGISTER_1_WR: out    vl_logic;
        oOTHER_REGISTER_1_NUM: out    vl_logic_vector(5 downto 0);
        iOTHER_REGISTER_1_FULL: in     vl_logic;
        iOTHER_REGISTER_1_COUNT: in     vl_logic_vector(2 downto 0);
        oNEXT_EX_BRANCH_VALID: out    vl_logic;
        oNEXT_EX_BRANCH_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_BRANCH_CMD: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_BRANCH_CC: out    vl_logic_vector(3 downto 0);
        oNEXT_EX_BRANCH_FLAG: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_BRANCH_SOURCE: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_PC     : out    vl_logic_vector(31 downto 0);
        iNEXT_EX_BRANCH_LOCK: in     vl_logic;
        iSCHE2_EX_BRANCH_VALID: in     vl_logic;
        iSCHE2_EX_BRANCH_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU1_VALID: out    vl_logic;
        oNEXT_EX_ALU1_WRITEBACK: out    vl_logic;
        oNEXT_EX_ALU1_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU1_CMD: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU1_AFE: out    vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU1_SYS_REG: out    vl_logic;
        oNEXT_EX_ALU1_LOGIC: out    vl_logic;
        oNEXT_EX_ALU1_SHIFT: out    vl_logic;
        oNEXT_EX_ALU1_ADDER: out    vl_logic;
        oNEXT_EX_ALU1_MUL: out    vl_logic;
        oNEXT_EX_ALU1_SDIV: out    vl_logic;
        oNEXT_EX_ALU1_UDIV: out    vl_logic;
        oNEXT_EX_ALU1_SOURCE0: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU1_SOURCE1: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU1_DESTINATION_SYSREG: out    vl_logic;
        oNEXT_EX_ALU1_LOGIC_DEST: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU1_DESTINATION_REGNAME: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU1_FLAGS_WRITEBACK: out    vl_logic;
        oNEXT_EX_ALU1_FLAGS_REGNAME: out    vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU1_PCR: out    vl_logic_vector(31 downto 0);
        iNEXT_EX_ALU1_LOCK: in     vl_logic;
        iSCHE2_EX_ALU1_VALID: in     vl_logic;
        iSCHE2_EX_ALU1_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iSCHE2_EX_ALU1_DESTINATION_SYSREG: in     vl_logic;
        iSCHE2_EX_ALU1_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iSCHE2_EX_ALU1_WRITEBACK: in     vl_logic;
        iSCHE2_EX_ALU1_DATA: in     vl_logic_vector(31 downto 0);
        iSCHE2_EX_ALU1_FLAG: in     vl_logic_vector(4 downto 0);
        iSCHE2_EX_ALU1_FLAGS_WRITEBACK: in     vl_logic;
        iSCHE2_EX_ALU1_FLAGS_REGNAME: in     vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU2_VALID: out    vl_logic;
        oNEXT_EX_ALU2_WRITEBACK: out    vl_logic;
        oNEXT_EX_ALU2_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU2_CMD: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU2_AFE: out    vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU2_SYS_REG: out    vl_logic;
        oNEXT_EX_ALU2_LOGIC: out    vl_logic;
        oNEXT_EX_ALU2_SHIFT: out    vl_logic;
        oNEXT_EX_ALU2_ADDER: out    vl_logic;
        oNEXT_EX_ALU2_SOURCE0: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU2_SOURCE1: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU2_DESTINATION_SYSREG: out    vl_logic;
        oNEXT_EX_ALU2_LOGIC_DEST: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU2_DESTINATION_REGNAME: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU2_FLAGS_WRITEBACK: out    vl_logic;
        oNEXT_EX_ALU2_FLAGS_REGNAME: out    vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU2_PCR: out    vl_logic_vector(31 downto 0);
        iNEXT_EX_ALU2_LOCK: in     vl_logic;
        iSCHE2_EX_ALU2_VALID: in     vl_logic;
        iSCHE2_EX_ALU2_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iSCHE2_EX_ALU2_DESTINATION_SYSREG: in     vl_logic;
        iSCHE2_EX_ALU2_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iSCHE2_EX_ALU2_WRITEBACK: in     vl_logic;
        iSCHE2_EX_ALU2_DATA: in     vl_logic_vector(31 downto 0);
        iSCHE2_EX_ALU2_FLAG: in     vl_logic_vector(4 downto 0);
        iSCHE2_EX_ALU2_FLAGS_WRITEBACK: in     vl_logic;
        iSCHE2_EX_ALU2_FLAGS_REGNAME: in     vl_logic_vector(3 downto 0);
        oNEXT_EX_ALU3_VALID: out    vl_logic;
        oNEXT_EX_ALU3_DESTINATION_SYSREG: out    vl_logic;
        oNEXT_EX_ALU3_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU3_CMD: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU3_SYS_LDST: out    vl_logic;
        oNEXT_EX_ALU3_LDST: out    vl_logic;
        oNEXT_EX_ALU3_SOURCE0: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU3_SOURCE1: out    vl_logic_vector(31 downto 0);
        oNEXT_EX_ALU3_ADV_ACTIVE: out    vl_logic;
        oNEXT_EX_ALU3_ADV_DATA: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU3_LOGIC_DEST: out    vl_logic_vector(4 downto 0);
        oNEXT_EX_ALU3_DESTINATION_REGNAME: out    vl_logic_vector(5 downto 0);
        oNEXT_EX_ALU3_PC: out    vl_logic_vector(31 downto 0);
        iNEXT_EX_ALU3_LOCK: in     vl_logic;
        iSCHE2_ALU3_VALID: in     vl_logic;
        iSCHE2_ALU3_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iSCHE2_ALU3_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iSCHE2_ALU3_DESTINATION_SYSREG: in     vl_logic;
        iSCHE2_ALU3_WRITEBACK: in     vl_logic;
        iSCHE2_ALU3_DATA: in     vl_logic_vector(31 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of CORE_ID : constant is 1;
end scheduler2;
