library verilog;
use verilog.vl_types.all;
entity \execute_port3_\ is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iRESET_SYNC     : in     vl_logic;
        iFREE_EX        : in     vl_logic;
        iFREE_SYSREG_NEW_SPR_VALID: in     vl_logic;
        iFREE_SYSREG_NEW_SPR: in     vl_logic_vector(31 downto 0);
        iSYSREG_TIDR    : in     vl_logic_vector(31 downto 0);
        iSYSREG_PSR     : in     vl_logic_vector(31 downto 0);
        iSYSREG_PDTR    : in     vl_logic_vector(31 downto 0);
        oSYSREG_SPR     : out    vl_logic_vector(31 downto 0);
        oDATAIO_REQ     : out    vl_logic;
        iDATAIO_BUSY    : in     vl_logic;
        oDATAIO_ORDER   : out    vl_logic_vector(1 downto 0);
        oDATAIO_MASK    : out    vl_logic_vector(3 downto 0);
        oDATAIO_RW      : out    vl_logic;
        oDATAIO_TID     : out    vl_logic_vector(13 downto 0);
        oDATAIO_MMUMOD  : out    vl_logic_vector(1 downto 0);
        oDATAIO_PDT     : out    vl_logic_vector(31 downto 0);
        oDATAIO_ADDR    : out    vl_logic_vector(31 downto 0);
        oDATAIO_DATA    : out    vl_logic_vector(31 downto 0);
        iDATAIO_REQ     : in     vl_logic;
        iDATAIO_DATA    : in     vl_logic_vector(31 downto 0);
        iPREVIOUS_EX_ALU3_VALID: in     vl_logic;
        iPREVIOUS_EX_ALU3_DESTINATION_SYSREG: in     vl_logic;
        iPREVIOUS_EX_ALU3_COMMIT_TAG: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_EX_ALU3_CMD: in     vl_logic_vector(4 downto 0);
        iPREVIOUS_EX_ALU3_SOURCE0: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_EX_ALU3_SOURCE1: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_EX_ALU3_ADV_ACTIVE: in     vl_logic;
        iPREVIOUS_EX_ALU3_ADV_DATA: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_EX_ALU3_DESTINATION_REGNAME: in     vl_logic_vector(5 downto 0);
        iPREVIOUS_EX_ALU3_PC: in     vl_logic_vector(31 downto 0);
        iPREVIOUS_EX_ALU3_SYS_LDST: in     vl_logic;
        iPREVIOUS_EX_ALU3_LDST: in     vl_logic;
        oPREVIOUS_EX_ALU3_LOCK: out    vl_logic;
        oSCHE1_ALU3_VALID: out    vl_logic;
        oSCHE1_ALU3_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oSCHE2_ALU3_VALID: out    vl_logic;
        oSCHE2_ALU3_COMMIT_TAG: out    vl_logic_vector(5 downto 0);
        oSCHE2_ALU3_DESTINATION_REGNAME: out    vl_logic_vector(5 downto 0);
        oSCHE2_ALU3_DESTINATION_SYSREG: out    vl_logic;
        oSCHE2_ALU3_WRITEBACK: out    vl_logic;
        oSCHE2_ALU3_DATA: out    vl_logic_vector(31 downto 0)
    );
end \execute_port3_\;
