library verilog;
use verilog.vl_types.all;
entity mimsr is
    port(
        iCLOCK          : in     vl_logic;
        inRESET         : in     vl_logic;
        iREQ_VALID      : in     vl_logic;
        oREQ_VALID      : out    vl_logic;
        oREQ_DATA       : out    vl_logic_vector(31 downto 0)
    );
end mimsr;
